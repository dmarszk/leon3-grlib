------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2015, Cobham Gaisler AB - all rights reserved.
--
-- ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN 
-- ACCORDANCE WITH THE GAISLER LICENSE AGREEMENT AND MUST BE APPROVED 
-- IN ADVANCE IN WRITING.
------------------------------------------------------------------------------


library ieee, cycloneiii;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use cycloneiii.cycloneiii_components.all;
library altera;
use altera.altera_primitives_components.all;

entity grlfpw_0_cycloneiii is
port(
  rst :  in std_logic;
  clk :  in std_logic;
  holdn :  in std_logic;
  cpi_flush :  in std_logic;
  cpi_exack :  in std_logic;
  cpi_a_rs1 : in std_logic_vector(4 downto 0);
  cpi_d_pc : in std_logic_vector(31 downto 0);
  cpi_d_inst : in std_logic_vector(31 downto 0);
  cpi_d_cnt : in std_logic_vector(1 downto 0);
  cpi_d_trap :  in std_logic;
  cpi_d_annul :  in std_logic;
  cpi_d_pv :  in std_logic;
  cpi_a_pc : in std_logic_vector(31 downto 0);
  cpi_a_inst : in std_logic_vector(31 downto 0);
  cpi_a_cnt : in std_logic_vector(1 downto 0);
  cpi_a_trap :  in std_logic;
  cpi_a_annul :  in std_logic;
  cpi_a_pv :  in std_logic;
  cpi_e_pc : in std_logic_vector(31 downto 0);
  cpi_e_inst : in std_logic_vector(31 downto 0);
  cpi_e_cnt : in std_logic_vector(1 downto 0);
  cpi_e_trap :  in std_logic;
  cpi_e_annul :  in std_logic;
  cpi_e_pv :  in std_logic;
  cpi_m_pc : in std_logic_vector(31 downto 0);
  cpi_m_inst : in std_logic_vector(31 downto 0);
  cpi_m_cnt : in std_logic_vector(1 downto 0);
  cpi_m_trap :  in std_logic;
  cpi_m_annul :  in std_logic;
  cpi_m_pv :  in std_logic;
  cpi_x_pc : in std_logic_vector(31 downto 0);
  cpi_x_inst : in std_logic_vector(31 downto 0);
  cpi_x_cnt : in std_logic_vector(1 downto 0);
  cpi_x_trap :  in std_logic;
  cpi_x_annul :  in std_logic;
  cpi_x_pv :  in std_logic;
  cpi_lddata : in std_logic_vector(31 downto 0);
  cpi_dbg_enable :  in std_logic;
  cpi_dbg_write :  in std_logic;
  cpi_dbg_fsr :  in std_logic;
  cpi_dbg_addr : in std_logic_vector(4 downto 0);
  cpi_dbg_data : in std_logic_vector(31 downto 0);
  cpo_data : out std_logic_vector(31 downto 0);
  cpo_exc :  out std_logic;
  cpo_cc : out std_logic_vector(1 downto 0);
  cpo_ccv :  out std_logic;
  cpo_ldlock :  out std_logic;
  cpo_holdn :  out std_logic;
  cpo_dbg_data : out std_logic_vector(31 downto 0);
  rfi1_rd1addr : out std_logic_vector(3 downto 0);
  rfi1_rd2addr : out std_logic_vector(3 downto 0);
  rfi1_wraddr : out std_logic_vector(3 downto 0);
  rfi1_wrdata : out std_logic_vector(31 downto 0);
  rfi1_ren1 :  out std_logic;
  rfi1_ren2 :  out std_logic;
  rfi1_wren :  out std_logic;
  rfi2_rd1addr : out std_logic_vector(3 downto 0);
  rfi2_rd2addr : out std_logic_vector(3 downto 0);
  rfi2_wraddr : out std_logic_vector(3 downto 0);
  rfi2_wrdata : out std_logic_vector(31 downto 0);
  rfi2_ren1 :  out std_logic;
  rfi2_ren2 :  out std_logic;
  rfi2_wren :  out std_logic;
  rfo1_data1 : in std_logic_vector(31 downto 0);
  rfo1_data2 : in std_logic_vector(31 downto 0);
  rfo2_data1 : in std_logic_vector(31 downto 0);
  rfo2_data2 : in std_logic_vector(31 downto 0));
end grlfpw_0_cycloneiii;

architecture beh of grlfpw_0_cycloneiii is
  signal devclrn : std_logic := '1';
  signal devpor : std_logic := '1';
  signal devoe : std_logic := '0';
  signal \GRLFPC20.FPI.OP2_X\ : std_logic_vector(63 downto 32);
  signal \GRLFPC20.R.FSR.RD\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.R.STATE\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.R.X.SEQERR\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.I.INST\ : std_logic_vector(31 downto 0);
  signal \GRLFPC20.R.FSR.TEM\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.I.EXC\ : std_logic_vector(5 downto 0);
  signal \GRLFPC20.R.FSR.AEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.A.RS1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.A.RS2\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.X.RDD\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.I.PC\ : std_logic_vector(31 downto 2);
  signal \GRLFPC20.R.FSR.CEXC\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.R.FSR.FTT\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.R.I.CC\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.R.I.RES\ : std_logic_vector(63 downto 0);
  signal \GRLFPC20.COMB.V.I.RES_6_X\ : std_logic_vector(63 to 63);
  signal \GRLFPC20.COMB.V.I.RES_1\ : std_logic_vector(63 to 63);
  signal \GRLFPC20.R.A.RF1REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC20.R.A.RF2REN\ : std_logic_vector(2 downto 1);
  signal \GRLFPC20.R.A.SEQERR\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.E.SEQERR\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.M.SEQERR\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.A.RDD\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.E.RDD\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.M.RDD\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.R.I.EXC_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.COMB.RS2_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.E.STDATA_1_0_X\ : std_logic_vector(31 downto 2);
  signal \GRLFPC20.COMB.V.E.STDATA_1_1\ : std_logic_vector(31 downto 2);
  signal \GRLFPC20.COMB.RS1_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.FSR.FCC_1\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.COMB.V.FSR.CEXC_1\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.FSR.CEXC_1_2\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\ : std_logic_vector(16 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\ : std_logic_vector(8 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\ : std_logic_vector(85 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\ : std_logic_vector(377 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\ : std_logic_vector(51 downto 30);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.MIXOIN\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_X\ : std_logic_vector(83 downto 81);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\ : std_logic_vector(80 downto 61);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\ : std_logic_vector(113 downto 61);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_V\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\ : std_logic_vector(12 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\ : std_logic_vector(12 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\ : std_logic_vector(257 downto 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.SUM_0_A2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.SUM\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\ : std_logic_vector(10 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\ : std_logic_vector(57 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_U\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_0_A2\ : std_logic_vector(19 to 19);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\ : std_logic_vector(257 downto 237);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\ : std_logic_vector(257 downto 250);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\ : std_logic_vector(83 downto 61);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.SUM_0_A2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0_A2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.COMB.V.A.RF1REN_1\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\ : std_logic_vector(8 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\ : std_logic_vector(56 downto 10);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\ : std_logic_vector(57 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\ : std_logic_vector(115 downto 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\ : std_logic_vector(115 downto 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\ : std_logic_vector(112 downto 58);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\ : std_logic_vector(55 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\ : std_logic_vector(54 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\ : std_logic_vector(22 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\ : std_logic_vector(57 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\ : std_logic_vector(57 downto 10);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\ : std_logic_vector(56 downto 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\ : std_logic_vector(55 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\ : std_logic_vector(55 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\ : std_logic_vector(68 to 68);
  signal \GRLFPC20.COMB.WRADDR_6_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.RS1_1_0_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.WRDATA_4_X\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.COMB.DBGDATA_4_0_X\ : std_logic_vector(31 downto 0);
  signal \GRLFPC20.WRDATA_0_X\ : std_logic_vector(63 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\ : std_logic_vector(57 downto 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\ : std_logic_vector(55 downto 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\ : std_logic_vector(62 downto 7);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\ : std_logic_vector(62 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\ : std_logic_vector(61 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\ : std_logic_vector(9 downto 3);
  signal \GRLFPC20.FPI.OP1_X\ : std_logic_vector(63 downto 32);
  signal \GRLFPC20.COMB.V.FSR.FCC_1_0_X\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.COMB.V.FSR.FCC_1_1_X\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.COMB.V.A.RF1REN_1_1_X\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.COMB.RF1REN_1_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.COMB.RF2REN_1_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.COMB.RF1REN_1_0_X\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.COMB.RF2REN_1_0_X\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STATUS\ : std_logic_vector(6 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT_0\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_27\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\ : std_logic_vector(9 downto 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\ : std_logic_vector(244 downto 115);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\ : std_logic_vector(257 downto 232);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\ : std_logic_vector(244 downto 237);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\ : std_logic_vector(8 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_0\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\ : std_logic_vector(9 downto 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2_1\ : std_logic_vector(9 to 9);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\ : std_logic_vector(9 downto 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\ : std_logic_vector(57 downto 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\ : std_logic_vector(2 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_18\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_21\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_25\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_15\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.NOTDIVC\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_3\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_6\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_9\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_14\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_12\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_0\ : std_logic_vector(12 to 12);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\ : std_logic_vector(4 to 4);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_0\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\ : std_logic_vector(2 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM_I\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19_U\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_0_A2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.QUOBITS\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\ : std_logic_vector(142 downto 141);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_V\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\ : std_logic_vector(59 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\ : std_logic_vector(58 downto 11);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\ : std_logic_vector(62 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\ : std_logic_vector(57 downto 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_0_A2\ : std_logic_vector(18 to 18);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\ : std_logic_vector(59 downto 12);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\ : std_logic_vector(62 downto 23);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_12\ : std_logic_vector(24 downto 23);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1_X\ : std_logic_vector(25 downto 23);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\ : std_logic_vector(57 downto 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_S\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0_D\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\ : std_logic_vector(67 to 67);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31_D\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0_D_0\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_15_D\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\ : std_logic_vector(8 downto 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31_S_0\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_4\ : std_logic_vector(6 downto 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_5\ : std_logic_vector(6 downto 5);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_0\ : std_logic_vector(4 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1\ : std_logic_vector(1 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_1\ : std_logic_vector(77 to 77);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_1\ : std_logic_vector(13 to 13);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV_0\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\ : std_logic_vector(56 to 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\ : std_logic_vector(75 to 75);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_0_A2\ : std_logic_vector(56 to 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\ : std_logic_vector(77 to 77);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_2_A\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\ : std_logic_vector(57 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\ : std_logic_vector(58 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\ : std_logic_vector(58 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\ : std_logic_vector(56 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\ : std_logic_vector(25 downto 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\ : std_logic_vector(54 downto 18);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_A\ : std_logic_vector(233 downto 113);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_A\ : std_logic_vector(48 downto 39);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\ : std_logic_vector(3 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_A\ : std_logic_vector(57 downto 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\ : std_logic_vector(32 downto 29);
  signal \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\ : std_logic_vector(4 downto 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_A\ : std_logic_vector(10 downto 8);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6_A\ : std_logic_vector(15 to 15);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1_A\ : std_logic_vector(1 to 1);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_A\ : std_logic_vector(0 to 0);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\ : std_logic_vector(54 downto 21);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\ : std_logic_vector(3 to 3);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_0_A\ : std_logic_vector(12 to 12);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4_A\ : std_logic_vector(56 to 56);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2_RETI\ : std_logic_vector(6 to 6);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\ : std_logic_vector(2 to 2);
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\ : std_logic_vector(78 to 78);
  signal CPO_DATAZ : std_logic_vector(31 downto 0);
  signal CPO_CCZ : std_logic_vector(1 downto 0);
  signal CPO_DBG_DATAZ : std_logic_vector(31 downto 0);
  signal RFI1_WRDATAZ : std_logic_vector(31 downto 0);
  signal RFI2_RD1ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_RD2ADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRADDRZ : std_logic_vector(3 downto 0);
  signal RFI2_WRDATAZ : std_logic_vector(31 downto 0);
  signal CLK_INTERNAL : std_logic ;
  signal CPI_FLUSH_INTERNAL : std_logic ;
  signal CPI_EXACK_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL : std_logic ;
  signal CPI_A_RS1_INTERNAL_0 : std_logic ;
  signal CPI_A_RS1_INTERNAL_1 : std_logic ;
  signal CPI_A_RS1_INTERNAL_2 : std_logic ;
  signal CPI_A_RS1_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL : std_logic ;
  signal CPI_D_PC_INTERNAL_0 : std_logic ;
  signal CPI_D_PC_INTERNAL_1 : std_logic ;
  signal CPI_D_PC_INTERNAL_2 : std_logic ;
  signal CPI_D_PC_INTERNAL_3 : std_logic ;
  signal CPI_D_PC_INTERNAL_4 : std_logic ;
  signal CPI_D_PC_INTERNAL_5 : std_logic ;
  signal CPI_D_PC_INTERNAL_6 : std_logic ;
  signal CPI_D_PC_INTERNAL_7 : std_logic ;
  signal CPI_D_PC_INTERNAL_8 : std_logic ;
  signal CPI_D_PC_INTERNAL_9 : std_logic ;
  signal CPI_D_PC_INTERNAL_10 : std_logic ;
  signal CPI_D_PC_INTERNAL_11 : std_logic ;
  signal CPI_D_PC_INTERNAL_12 : std_logic ;
  signal CPI_D_PC_INTERNAL_13 : std_logic ;
  signal CPI_D_PC_INTERNAL_14 : std_logic ;
  signal CPI_D_PC_INTERNAL_15 : std_logic ;
  signal CPI_D_PC_INTERNAL_16 : std_logic ;
  signal CPI_D_PC_INTERNAL_17 : std_logic ;
  signal CPI_D_PC_INTERNAL_18 : std_logic ;
  signal CPI_D_PC_INTERNAL_19 : std_logic ;
  signal CPI_D_PC_INTERNAL_20 : std_logic ;
  signal CPI_D_PC_INTERNAL_21 : std_logic ;
  signal CPI_D_PC_INTERNAL_22 : std_logic ;
  signal CPI_D_PC_INTERNAL_23 : std_logic ;
  signal CPI_D_PC_INTERNAL_24 : std_logic ;
  signal CPI_D_PC_INTERNAL_25 : std_logic ;
  signal CPI_D_PC_INTERNAL_26 : std_logic ;
  signal CPI_D_PC_INTERNAL_27 : std_logic ;
  signal CPI_D_PC_INTERNAL_28 : std_logic ;
  signal CPI_D_PC_INTERNAL_29 : std_logic ;
  signal CPI_D_PC_INTERNAL_30 : std_logic ;
  signal CPI_D_INST_INTERNAL : std_logic ;
  signal CPI_D_INST_INTERNAL_0 : std_logic ;
  signal CPI_D_INST_INTERNAL_1 : std_logic ;
  signal CPI_D_INST_INTERNAL_2 : std_logic ;
  signal CPI_D_INST_INTERNAL_3 : std_logic ;
  signal CPI_D_INST_INTERNAL_4 : std_logic ;
  signal CPI_D_INST_INTERNAL_5 : std_logic ;
  signal CPI_D_INST_INTERNAL_6 : std_logic ;
  signal CPI_D_INST_INTERNAL_7 : std_logic ;
  signal CPI_D_INST_INTERNAL_8 : std_logic ;
  signal CPI_D_INST_INTERNAL_9 : std_logic ;
  signal CPI_D_INST_INTERNAL_10 : std_logic ;
  signal CPI_D_INST_INTERNAL_11 : std_logic ;
  signal CPI_D_INST_INTERNAL_12 : std_logic ;
  signal CPI_D_INST_INTERNAL_13 : std_logic ;
  signal CPI_D_INST_INTERNAL_14 : std_logic ;
  signal CPI_D_INST_INTERNAL_15 : std_logic ;
  signal CPI_D_INST_INTERNAL_16 : std_logic ;
  signal CPI_D_INST_INTERNAL_17 : std_logic ;
  signal CPI_D_INST_INTERNAL_18 : std_logic ;
  signal CPI_D_INST_INTERNAL_19 : std_logic ;
  signal CPI_D_INST_INTERNAL_20 : std_logic ;
  signal CPI_D_INST_INTERNAL_21 : std_logic ;
  signal CPI_D_INST_INTERNAL_22 : std_logic ;
  signal CPI_D_INST_INTERNAL_23 : std_logic ;
  signal CPI_D_INST_INTERNAL_24 : std_logic ;
  signal CPI_D_INST_INTERNAL_25 : std_logic ;
  signal CPI_D_INST_INTERNAL_26 : std_logic ;
  signal CPI_D_INST_INTERNAL_27 : std_logic ;
  signal CPI_D_INST_INTERNAL_28 : std_logic ;
  signal CPI_D_INST_INTERNAL_29 : std_logic ;
  signal CPI_D_INST_INTERNAL_30 : std_logic ;
  signal CPI_D_CNT_INTERNAL : std_logic ;
  signal CPI_D_CNT_INTERNAL_0 : std_logic ;
  signal CPI_D_TRAP_INTERNAL : std_logic ;
  signal CPI_D_ANNUL_INTERNAL : std_logic ;
  signal CPI_D_PV_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL : std_logic ;
  signal CPI_A_PC_INTERNAL_0 : std_logic ;
  signal CPI_A_PC_INTERNAL_1 : std_logic ;
  signal CPI_A_PC_INTERNAL_2 : std_logic ;
  signal CPI_A_PC_INTERNAL_3 : std_logic ;
  signal CPI_A_PC_INTERNAL_4 : std_logic ;
  signal CPI_A_PC_INTERNAL_5 : std_logic ;
  signal CPI_A_PC_INTERNAL_6 : std_logic ;
  signal CPI_A_PC_INTERNAL_7 : std_logic ;
  signal CPI_A_PC_INTERNAL_8 : std_logic ;
  signal CPI_A_PC_INTERNAL_9 : std_logic ;
  signal CPI_A_PC_INTERNAL_10 : std_logic ;
  signal CPI_A_PC_INTERNAL_11 : std_logic ;
  signal CPI_A_PC_INTERNAL_12 : std_logic ;
  signal CPI_A_PC_INTERNAL_13 : std_logic ;
  signal CPI_A_PC_INTERNAL_14 : std_logic ;
  signal CPI_A_PC_INTERNAL_15 : std_logic ;
  signal CPI_A_PC_INTERNAL_16 : std_logic ;
  signal CPI_A_PC_INTERNAL_17 : std_logic ;
  signal CPI_A_PC_INTERNAL_18 : std_logic ;
  signal CPI_A_PC_INTERNAL_19 : std_logic ;
  signal CPI_A_PC_INTERNAL_20 : std_logic ;
  signal CPI_A_PC_INTERNAL_21 : std_logic ;
  signal CPI_A_PC_INTERNAL_22 : std_logic ;
  signal CPI_A_PC_INTERNAL_23 : std_logic ;
  signal CPI_A_PC_INTERNAL_24 : std_logic ;
  signal CPI_A_PC_INTERNAL_25 : std_logic ;
  signal CPI_A_PC_INTERNAL_26 : std_logic ;
  signal CPI_A_PC_INTERNAL_27 : std_logic ;
  signal CPI_A_PC_INTERNAL_28 : std_logic ;
  signal CPI_A_PC_INTERNAL_29 : std_logic ;
  signal CPI_A_PC_INTERNAL_30 : std_logic ;
  signal CPI_A_INST_INTERNAL : std_logic ;
  signal CPI_A_INST_INTERNAL_0 : std_logic ;
  signal CPI_A_INST_INTERNAL_1 : std_logic ;
  signal CPI_A_INST_INTERNAL_2 : std_logic ;
  signal CPI_A_INST_INTERNAL_3 : std_logic ;
  signal CPI_A_INST_INTERNAL_4 : std_logic ;
  signal CPI_A_INST_INTERNAL_5 : std_logic ;
  signal CPI_A_INST_INTERNAL_6 : std_logic ;
  signal CPI_A_INST_INTERNAL_7 : std_logic ;
  signal CPI_A_INST_INTERNAL_8 : std_logic ;
  signal CPI_A_INST_INTERNAL_9 : std_logic ;
  signal CPI_A_INST_INTERNAL_10 : std_logic ;
  signal CPI_A_INST_INTERNAL_11 : std_logic ;
  signal CPI_A_INST_INTERNAL_12 : std_logic ;
  signal CPI_A_INST_INTERNAL_13 : std_logic ;
  signal CPI_A_INST_INTERNAL_14 : std_logic ;
  signal CPI_A_INST_INTERNAL_15 : std_logic ;
  signal CPI_A_INST_INTERNAL_16 : std_logic ;
  signal CPI_A_INST_INTERNAL_17 : std_logic ;
  signal CPI_A_INST_INTERNAL_18 : std_logic ;
  signal CPI_A_INST_INTERNAL_19 : std_logic ;
  signal CPI_A_INST_INTERNAL_20 : std_logic ;
  signal CPI_A_INST_INTERNAL_21 : std_logic ;
  signal CPI_A_INST_INTERNAL_22 : std_logic ;
  signal CPI_A_INST_INTERNAL_23 : std_logic ;
  signal CPI_A_INST_INTERNAL_24 : std_logic ;
  signal CPI_A_INST_INTERNAL_25 : std_logic ;
  signal CPI_A_INST_INTERNAL_26 : std_logic ;
  signal CPI_A_INST_INTERNAL_27 : std_logic ;
  signal CPI_A_INST_INTERNAL_28 : std_logic ;
  signal CPI_A_INST_INTERNAL_29 : std_logic ;
  signal CPI_A_INST_INTERNAL_30 : std_logic ;
  signal CPI_A_CNT_INTERNAL : std_logic ;
  signal CPI_A_CNT_INTERNAL_0 : std_logic ;
  signal CPI_A_TRAP_INTERNAL : std_logic ;
  signal CPI_A_ANNUL_INTERNAL : std_logic ;
  signal CPI_A_PV_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL : std_logic ;
  signal CPI_E_PC_INTERNAL_0 : std_logic ;
  signal CPI_E_PC_INTERNAL_1 : std_logic ;
  signal CPI_E_PC_INTERNAL_2 : std_logic ;
  signal CPI_E_PC_INTERNAL_3 : std_logic ;
  signal CPI_E_PC_INTERNAL_4 : std_logic ;
  signal CPI_E_PC_INTERNAL_5 : std_logic ;
  signal CPI_E_PC_INTERNAL_6 : std_logic ;
  signal CPI_E_PC_INTERNAL_7 : std_logic ;
  signal CPI_E_PC_INTERNAL_8 : std_logic ;
  signal CPI_E_PC_INTERNAL_9 : std_logic ;
  signal CPI_E_PC_INTERNAL_10 : std_logic ;
  signal CPI_E_PC_INTERNAL_11 : std_logic ;
  signal CPI_E_PC_INTERNAL_12 : std_logic ;
  signal CPI_E_PC_INTERNAL_13 : std_logic ;
  signal CPI_E_PC_INTERNAL_14 : std_logic ;
  signal CPI_E_PC_INTERNAL_15 : std_logic ;
  signal CPI_E_PC_INTERNAL_16 : std_logic ;
  signal CPI_E_PC_INTERNAL_17 : std_logic ;
  signal CPI_E_PC_INTERNAL_18 : std_logic ;
  signal CPI_E_PC_INTERNAL_19 : std_logic ;
  signal CPI_E_PC_INTERNAL_20 : std_logic ;
  signal CPI_E_PC_INTERNAL_21 : std_logic ;
  signal CPI_E_PC_INTERNAL_22 : std_logic ;
  signal CPI_E_PC_INTERNAL_23 : std_logic ;
  signal CPI_E_PC_INTERNAL_24 : std_logic ;
  signal CPI_E_PC_INTERNAL_25 : std_logic ;
  signal CPI_E_PC_INTERNAL_26 : std_logic ;
  signal CPI_E_PC_INTERNAL_27 : std_logic ;
  signal CPI_E_PC_INTERNAL_28 : std_logic ;
  signal CPI_E_PC_INTERNAL_29 : std_logic ;
  signal CPI_E_PC_INTERNAL_30 : std_logic ;
  signal CPI_E_INST_INTERNAL : std_logic ;
  signal CPI_E_INST_INTERNAL_0 : std_logic ;
  signal CPI_E_INST_INTERNAL_1 : std_logic ;
  signal CPI_E_INST_INTERNAL_2 : std_logic ;
  signal CPI_E_INST_INTERNAL_3 : std_logic ;
  signal CPI_E_INST_INTERNAL_4 : std_logic ;
  signal CPI_E_INST_INTERNAL_5 : std_logic ;
  signal CPI_E_INST_INTERNAL_6 : std_logic ;
  signal CPI_E_INST_INTERNAL_7 : std_logic ;
  signal CPI_E_INST_INTERNAL_8 : std_logic ;
  signal CPI_E_INST_INTERNAL_9 : std_logic ;
  signal CPI_E_INST_INTERNAL_10 : std_logic ;
  signal CPI_E_INST_INTERNAL_11 : std_logic ;
  signal CPI_E_INST_INTERNAL_12 : std_logic ;
  signal CPI_E_INST_INTERNAL_13 : std_logic ;
  signal CPI_E_INST_INTERNAL_14 : std_logic ;
  signal CPI_E_INST_INTERNAL_15 : std_logic ;
  signal CPI_E_INST_INTERNAL_16 : std_logic ;
  signal CPI_E_INST_INTERNAL_17 : std_logic ;
  signal CPI_E_INST_INTERNAL_18 : std_logic ;
  signal CPI_E_INST_INTERNAL_19 : std_logic ;
  signal CPI_E_INST_INTERNAL_20 : std_logic ;
  signal CPI_E_INST_INTERNAL_21 : std_logic ;
  signal CPI_E_INST_INTERNAL_22 : std_logic ;
  signal CPI_E_INST_INTERNAL_23 : std_logic ;
  signal CPI_E_INST_INTERNAL_24 : std_logic ;
  signal CPI_E_INST_INTERNAL_25 : std_logic ;
  signal CPI_E_INST_INTERNAL_26 : std_logic ;
  signal CPI_E_INST_INTERNAL_27 : std_logic ;
  signal CPI_E_INST_INTERNAL_28 : std_logic ;
  signal CPI_E_INST_INTERNAL_29 : std_logic ;
  signal CPI_E_INST_INTERNAL_30 : std_logic ;
  signal CPI_E_CNT_INTERNAL : std_logic ;
  signal CPI_E_CNT_INTERNAL_0 : std_logic ;
  signal CPI_E_TRAP_INTERNAL : std_logic ;
  signal CPI_E_ANNUL_INTERNAL : std_logic ;
  signal CPI_E_PV_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL : std_logic ;
  signal CPI_M_PC_INTERNAL_0 : std_logic ;
  signal CPI_M_PC_INTERNAL_1 : std_logic ;
  signal CPI_M_PC_INTERNAL_2 : std_logic ;
  signal CPI_M_PC_INTERNAL_3 : std_logic ;
  signal CPI_M_PC_INTERNAL_4 : std_logic ;
  signal CPI_M_PC_INTERNAL_5 : std_logic ;
  signal CPI_M_PC_INTERNAL_6 : std_logic ;
  signal CPI_M_PC_INTERNAL_7 : std_logic ;
  signal CPI_M_PC_INTERNAL_8 : std_logic ;
  signal CPI_M_PC_INTERNAL_9 : std_logic ;
  signal CPI_M_PC_INTERNAL_10 : std_logic ;
  signal CPI_M_PC_INTERNAL_11 : std_logic ;
  signal CPI_M_PC_INTERNAL_12 : std_logic ;
  signal CPI_M_PC_INTERNAL_13 : std_logic ;
  signal CPI_M_PC_INTERNAL_14 : std_logic ;
  signal CPI_M_PC_INTERNAL_15 : std_logic ;
  signal CPI_M_PC_INTERNAL_16 : std_logic ;
  signal CPI_M_PC_INTERNAL_17 : std_logic ;
  signal CPI_M_PC_INTERNAL_18 : std_logic ;
  signal CPI_M_PC_INTERNAL_19 : std_logic ;
  signal CPI_M_PC_INTERNAL_20 : std_logic ;
  signal CPI_M_PC_INTERNAL_21 : std_logic ;
  signal CPI_M_PC_INTERNAL_22 : std_logic ;
  signal CPI_M_PC_INTERNAL_23 : std_logic ;
  signal CPI_M_PC_INTERNAL_24 : std_logic ;
  signal CPI_M_PC_INTERNAL_25 : std_logic ;
  signal CPI_M_PC_INTERNAL_26 : std_logic ;
  signal CPI_M_PC_INTERNAL_27 : std_logic ;
  signal CPI_M_PC_INTERNAL_28 : std_logic ;
  signal CPI_M_PC_INTERNAL_29 : std_logic ;
  signal CPI_M_PC_INTERNAL_30 : std_logic ;
  signal CPI_M_INST_INTERNAL : std_logic ;
  signal CPI_M_INST_INTERNAL_0 : std_logic ;
  signal CPI_M_INST_INTERNAL_1 : std_logic ;
  signal CPI_M_INST_INTERNAL_2 : std_logic ;
  signal CPI_M_INST_INTERNAL_3 : std_logic ;
  signal CPI_M_INST_INTERNAL_4 : std_logic ;
  signal CPI_M_INST_INTERNAL_5 : std_logic ;
  signal CPI_M_INST_INTERNAL_6 : std_logic ;
  signal CPI_M_INST_INTERNAL_7 : std_logic ;
  signal CPI_M_INST_INTERNAL_8 : std_logic ;
  signal CPI_M_INST_INTERNAL_9 : std_logic ;
  signal CPI_M_INST_INTERNAL_10 : std_logic ;
  signal CPI_M_INST_INTERNAL_11 : std_logic ;
  signal CPI_M_INST_INTERNAL_12 : std_logic ;
  signal CPI_M_INST_INTERNAL_13 : std_logic ;
  signal CPI_M_INST_INTERNAL_14 : std_logic ;
  signal CPI_M_INST_INTERNAL_15 : std_logic ;
  signal CPI_M_INST_INTERNAL_16 : std_logic ;
  signal CPI_M_INST_INTERNAL_17 : std_logic ;
  signal CPI_M_INST_INTERNAL_18 : std_logic ;
  signal CPI_M_INST_INTERNAL_19 : std_logic ;
  signal CPI_M_INST_INTERNAL_20 : std_logic ;
  signal CPI_M_INST_INTERNAL_21 : std_logic ;
  signal CPI_M_INST_INTERNAL_22 : std_logic ;
  signal CPI_M_INST_INTERNAL_23 : std_logic ;
  signal CPI_M_INST_INTERNAL_24 : std_logic ;
  signal CPI_M_INST_INTERNAL_25 : std_logic ;
  signal CPI_M_INST_INTERNAL_26 : std_logic ;
  signal CPI_M_INST_INTERNAL_27 : std_logic ;
  signal CPI_M_INST_INTERNAL_28 : std_logic ;
  signal CPI_M_INST_INTERNAL_29 : std_logic ;
  signal CPI_M_INST_INTERNAL_30 : std_logic ;
  signal CPI_M_CNT_INTERNAL : std_logic ;
  signal CPI_M_CNT_INTERNAL_0 : std_logic ;
  signal CPI_M_TRAP_INTERNAL : std_logic ;
  signal CPI_M_ANNUL_INTERNAL : std_logic ;
  signal CPI_M_PV_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL : std_logic ;
  signal CPI_X_PC_INTERNAL_0 : std_logic ;
  signal CPI_X_PC_INTERNAL_1 : std_logic ;
  signal CPI_X_PC_INTERNAL_2 : std_logic ;
  signal CPI_X_PC_INTERNAL_3 : std_logic ;
  signal CPI_X_PC_INTERNAL_4 : std_logic ;
  signal CPI_X_PC_INTERNAL_5 : std_logic ;
  signal CPI_X_PC_INTERNAL_6 : std_logic ;
  signal CPI_X_PC_INTERNAL_7 : std_logic ;
  signal CPI_X_PC_INTERNAL_8 : std_logic ;
  signal CPI_X_PC_INTERNAL_9 : std_logic ;
  signal CPI_X_PC_INTERNAL_10 : std_logic ;
  signal CPI_X_PC_INTERNAL_11 : std_logic ;
  signal CPI_X_PC_INTERNAL_12 : std_logic ;
  signal CPI_X_PC_INTERNAL_13 : std_logic ;
  signal CPI_X_PC_INTERNAL_14 : std_logic ;
  signal CPI_X_PC_INTERNAL_15 : std_logic ;
  signal CPI_X_PC_INTERNAL_16 : std_logic ;
  signal CPI_X_PC_INTERNAL_17 : std_logic ;
  signal CPI_X_PC_INTERNAL_18 : std_logic ;
  signal CPI_X_PC_INTERNAL_19 : std_logic ;
  signal CPI_X_PC_INTERNAL_20 : std_logic ;
  signal CPI_X_PC_INTERNAL_21 : std_logic ;
  signal CPI_X_PC_INTERNAL_22 : std_logic ;
  signal CPI_X_PC_INTERNAL_23 : std_logic ;
  signal CPI_X_PC_INTERNAL_24 : std_logic ;
  signal CPI_X_PC_INTERNAL_25 : std_logic ;
  signal CPI_X_PC_INTERNAL_26 : std_logic ;
  signal CPI_X_PC_INTERNAL_27 : std_logic ;
  signal CPI_X_PC_INTERNAL_28 : std_logic ;
  signal CPI_X_PC_INTERNAL_29 : std_logic ;
  signal CPI_X_PC_INTERNAL_30 : std_logic ;
  signal CPI_X_INST_INTERNAL : std_logic ;
  signal CPI_X_INST_INTERNAL_0 : std_logic ;
  signal CPI_X_INST_INTERNAL_1 : std_logic ;
  signal CPI_X_INST_INTERNAL_2 : std_logic ;
  signal CPI_X_INST_INTERNAL_3 : std_logic ;
  signal CPI_X_INST_INTERNAL_4 : std_logic ;
  signal CPI_X_INST_INTERNAL_5 : std_logic ;
  signal CPI_X_INST_INTERNAL_6 : std_logic ;
  signal CPI_X_INST_INTERNAL_7 : std_logic ;
  signal CPI_X_INST_INTERNAL_8 : std_logic ;
  signal CPI_X_INST_INTERNAL_9 : std_logic ;
  signal CPI_X_INST_INTERNAL_10 : std_logic ;
  signal CPI_X_INST_INTERNAL_11 : std_logic ;
  signal CPI_X_INST_INTERNAL_12 : std_logic ;
  signal CPI_X_INST_INTERNAL_13 : std_logic ;
  signal CPI_X_INST_INTERNAL_14 : std_logic ;
  signal CPI_X_INST_INTERNAL_15 : std_logic ;
  signal CPI_X_INST_INTERNAL_16 : std_logic ;
  signal CPI_X_INST_INTERNAL_17 : std_logic ;
  signal CPI_X_INST_INTERNAL_18 : std_logic ;
  signal CPI_X_INST_INTERNAL_19 : std_logic ;
  signal CPI_X_INST_INTERNAL_20 : std_logic ;
  signal CPI_X_INST_INTERNAL_21 : std_logic ;
  signal CPI_X_INST_INTERNAL_22 : std_logic ;
  signal CPI_X_INST_INTERNAL_23 : std_logic ;
  signal CPI_X_INST_INTERNAL_24 : std_logic ;
  signal CPI_X_INST_INTERNAL_25 : std_logic ;
  signal CPI_X_INST_INTERNAL_26 : std_logic ;
  signal CPI_X_INST_INTERNAL_27 : std_logic ;
  signal CPI_X_INST_INTERNAL_28 : std_logic ;
  signal CPI_X_INST_INTERNAL_29 : std_logic ;
  signal CPI_X_INST_INTERNAL_30 : std_logic ;
  signal CPI_X_CNT_INTERNAL : std_logic ;
  signal CPI_X_CNT_INTERNAL_0 : std_logic ;
  signal CPI_X_TRAP_INTERNAL : std_logic ;
  signal CPI_X_ANNUL_INTERNAL : std_logic ;
  signal CPI_X_PV_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL : std_logic ;
  signal CPI_LDDATA_INTERNAL_0 : std_logic ;
  signal CPI_LDDATA_INTERNAL_1 : std_logic ;
  signal CPI_LDDATA_INTERNAL_2 : std_logic ;
  signal CPI_LDDATA_INTERNAL_3 : std_logic ;
  signal CPI_LDDATA_INTERNAL_4 : std_logic ;
  signal CPI_LDDATA_INTERNAL_5 : std_logic ;
  signal CPI_LDDATA_INTERNAL_6 : std_logic ;
  signal CPI_LDDATA_INTERNAL_7 : std_logic ;
  signal CPI_LDDATA_INTERNAL_8 : std_logic ;
  signal CPI_LDDATA_INTERNAL_9 : std_logic ;
  signal CPI_LDDATA_INTERNAL_10 : std_logic ;
  signal CPI_LDDATA_INTERNAL_11 : std_logic ;
  signal CPI_LDDATA_INTERNAL_12 : std_logic ;
  signal CPI_LDDATA_INTERNAL_13 : std_logic ;
  signal CPI_LDDATA_INTERNAL_14 : std_logic ;
  signal CPI_LDDATA_INTERNAL_15 : std_logic ;
  signal CPI_LDDATA_INTERNAL_16 : std_logic ;
  signal CPI_LDDATA_INTERNAL_17 : std_logic ;
  signal CPI_LDDATA_INTERNAL_18 : std_logic ;
  signal CPI_LDDATA_INTERNAL_19 : std_logic ;
  signal CPI_LDDATA_INTERNAL_20 : std_logic ;
  signal CPI_LDDATA_INTERNAL_21 : std_logic ;
  signal CPI_LDDATA_INTERNAL_22 : std_logic ;
  signal CPI_LDDATA_INTERNAL_23 : std_logic ;
  signal CPI_LDDATA_INTERNAL_24 : std_logic ;
  signal CPI_LDDATA_INTERNAL_25 : std_logic ;
  signal CPI_LDDATA_INTERNAL_26 : std_logic ;
  signal CPI_LDDATA_INTERNAL_27 : std_logic ;
  signal CPI_LDDATA_INTERNAL_28 : std_logic ;
  signal CPI_LDDATA_INTERNAL_29 : std_logic ;
  signal CPI_LDDATA_INTERNAL_30 : std_logic ;
  signal CPI_DBG_ENABLE_INTERNAL : std_logic ;
  signal CPI_DBG_WRITE_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_0 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_1 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_2 : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_0 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_1 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_2 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_3 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_4 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_5 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_6 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_7 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_8 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_9 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_10 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_11 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_12 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_13 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_14 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_15 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_16 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_17 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_18 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_19 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_20 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_21 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_22 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_23 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_24 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_25 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_26 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_27 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_28 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_29 : std_logic ;
  signal CPI_DBG_DATA_INTERNAL_30 : std_logic ;
  signal RFO1_DATA1_INTERNAL : std_logic ;
  signal RFO1_DATA1_INTERNAL_0 : std_logic ;
  signal RFO1_DATA1_INTERNAL_1 : std_logic ;
  signal RFO1_DATA1_INTERNAL_2 : std_logic ;
  signal RFO1_DATA1_INTERNAL_3 : std_logic ;
  signal RFO1_DATA1_INTERNAL_4 : std_logic ;
  signal RFO1_DATA1_INTERNAL_5 : std_logic ;
  signal RFO1_DATA1_INTERNAL_6 : std_logic ;
  signal RFO1_DATA1_INTERNAL_7 : std_logic ;
  signal RFO1_DATA1_INTERNAL_8 : std_logic ;
  signal RFO1_DATA1_INTERNAL_9 : std_logic ;
  signal RFO1_DATA1_INTERNAL_10 : std_logic ;
  signal RFO1_DATA1_INTERNAL_11 : std_logic ;
  signal RFO1_DATA1_INTERNAL_12 : std_logic ;
  signal RFO1_DATA1_INTERNAL_13 : std_logic ;
  signal RFO1_DATA1_INTERNAL_14 : std_logic ;
  signal RFO1_DATA1_INTERNAL_15 : std_logic ;
  signal RFO1_DATA1_INTERNAL_16 : std_logic ;
  signal RFO1_DATA1_INTERNAL_17 : std_logic ;
  signal RFO1_DATA1_INTERNAL_18 : std_logic ;
  signal RFO1_DATA1_INTERNAL_19 : std_logic ;
  signal RFO1_DATA1_INTERNAL_20 : std_logic ;
  signal RFO1_DATA1_INTERNAL_21 : std_logic ;
  signal RFO1_DATA1_INTERNAL_22 : std_logic ;
  signal RFO1_DATA1_INTERNAL_23 : std_logic ;
  signal RFO1_DATA1_INTERNAL_24 : std_logic ;
  signal RFO1_DATA1_INTERNAL_25 : std_logic ;
  signal RFO1_DATA1_INTERNAL_26 : std_logic ;
  signal RFO1_DATA1_INTERNAL_27 : std_logic ;
  signal RFO1_DATA1_INTERNAL_28 : std_logic ;
  signal RFO1_DATA1_INTERNAL_29 : std_logic ;
  signal RFO1_DATA1_INTERNAL_30 : std_logic ;
  signal RFO1_DATA2_INTERNAL : std_logic ;
  signal RFO1_DATA2_INTERNAL_0 : std_logic ;
  signal RFO1_DATA2_INTERNAL_1 : std_logic ;
  signal RFO1_DATA2_INTERNAL_2 : std_logic ;
  signal RFO1_DATA2_INTERNAL_3 : std_logic ;
  signal RFO1_DATA2_INTERNAL_4 : std_logic ;
  signal RFO1_DATA2_INTERNAL_5 : std_logic ;
  signal RFO1_DATA2_INTERNAL_6 : std_logic ;
  signal RFO1_DATA2_INTERNAL_7 : std_logic ;
  signal RFO1_DATA2_INTERNAL_8 : std_logic ;
  signal RFO1_DATA2_INTERNAL_9 : std_logic ;
  signal RFO1_DATA2_INTERNAL_10 : std_logic ;
  signal RFO1_DATA2_INTERNAL_11 : std_logic ;
  signal RFO1_DATA2_INTERNAL_12 : std_logic ;
  signal RFO1_DATA2_INTERNAL_13 : std_logic ;
  signal RFO1_DATA2_INTERNAL_14 : std_logic ;
  signal RFO1_DATA2_INTERNAL_15 : std_logic ;
  signal RFO1_DATA2_INTERNAL_16 : std_logic ;
  signal RFO1_DATA2_INTERNAL_17 : std_logic ;
  signal RFO1_DATA2_INTERNAL_18 : std_logic ;
  signal RFO1_DATA2_INTERNAL_19 : std_logic ;
  signal RFO1_DATA2_INTERNAL_20 : std_logic ;
  signal RFO1_DATA2_INTERNAL_21 : std_logic ;
  signal RFO1_DATA2_INTERNAL_22 : std_logic ;
  signal RFO1_DATA2_INTERNAL_23 : std_logic ;
  signal RFO1_DATA2_INTERNAL_24 : std_logic ;
  signal RFO1_DATA2_INTERNAL_25 : std_logic ;
  signal RFO1_DATA2_INTERNAL_26 : std_logic ;
  signal RFO1_DATA2_INTERNAL_27 : std_logic ;
  signal RFO1_DATA2_INTERNAL_28 : std_logic ;
  signal RFO1_DATA2_INTERNAL_29 : std_logic ;
  signal RFO1_DATA2_INTERNAL_30 : std_logic ;
  signal RFO2_DATA1_INTERNAL : std_logic ;
  signal RFO2_DATA1_INTERNAL_0 : std_logic ;
  signal RFO2_DATA1_INTERNAL_1 : std_logic ;
  signal RFO2_DATA1_INTERNAL_2 : std_logic ;
  signal RFO2_DATA1_INTERNAL_3 : std_logic ;
  signal RFO2_DATA1_INTERNAL_4 : std_logic ;
  signal RFO2_DATA1_INTERNAL_5 : std_logic ;
  signal RFO2_DATA1_INTERNAL_6 : std_logic ;
  signal RFO2_DATA1_INTERNAL_7 : std_logic ;
  signal RFO2_DATA1_INTERNAL_8 : std_logic ;
  signal RFO2_DATA1_INTERNAL_9 : std_logic ;
  signal RFO2_DATA1_INTERNAL_10 : std_logic ;
  signal RFO2_DATA1_INTERNAL_11 : std_logic ;
  signal RFO2_DATA1_INTERNAL_12 : std_logic ;
  signal RFO2_DATA1_INTERNAL_13 : std_logic ;
  signal RFO2_DATA1_INTERNAL_14 : std_logic ;
  signal RFO2_DATA1_INTERNAL_15 : std_logic ;
  signal RFO2_DATA1_INTERNAL_16 : std_logic ;
  signal RFO2_DATA1_INTERNAL_17 : std_logic ;
  signal RFO2_DATA1_INTERNAL_18 : std_logic ;
  signal RFO2_DATA1_INTERNAL_19 : std_logic ;
  signal RFO2_DATA1_INTERNAL_20 : std_logic ;
  signal RFO2_DATA1_INTERNAL_21 : std_logic ;
  signal RFO2_DATA1_INTERNAL_22 : std_logic ;
  signal RFO2_DATA1_INTERNAL_23 : std_logic ;
  signal RFO2_DATA1_INTERNAL_24 : std_logic ;
  signal RFO2_DATA1_INTERNAL_25 : std_logic ;
  signal RFO2_DATA1_INTERNAL_26 : std_logic ;
  signal RFO2_DATA1_INTERNAL_27 : std_logic ;
  signal RFO2_DATA1_INTERNAL_28 : std_logic ;
  signal RFO2_DATA1_INTERNAL_29 : std_logic ;
  signal RFO2_DATA1_INTERNAL_30 : std_logic ;
  signal RFO2_DATA2_INTERNAL : std_logic ;
  signal RFO2_DATA2_INTERNAL_0 : std_logic ;
  signal RFO2_DATA2_INTERNAL_1 : std_logic ;
  signal RFO2_DATA2_INTERNAL_2 : std_logic ;
  signal RFO2_DATA2_INTERNAL_3 : std_logic ;
  signal RFO2_DATA2_INTERNAL_4 : std_logic ;
  signal RFO2_DATA2_INTERNAL_5 : std_logic ;
  signal RFO2_DATA2_INTERNAL_6 : std_logic ;
  signal RFO2_DATA2_INTERNAL_7 : std_logic ;
  signal RFO2_DATA2_INTERNAL_8 : std_logic ;
  signal RFO2_DATA2_INTERNAL_9 : std_logic ;
  signal RFO2_DATA2_INTERNAL_10 : std_logic ;
  signal RFO2_DATA2_INTERNAL_11 : std_logic ;
  signal RFO2_DATA2_INTERNAL_12 : std_logic ;
  signal RFO2_DATA2_INTERNAL_13 : std_logic ;
  signal RFO2_DATA2_INTERNAL_14 : std_logic ;
  signal RFO2_DATA2_INTERNAL_15 : std_logic ;
  signal RFO2_DATA2_INTERNAL_16 : std_logic ;
  signal RFO2_DATA2_INTERNAL_17 : std_logic ;
  signal RFO2_DATA2_INTERNAL_18 : std_logic ;
  signal RFO2_DATA2_INTERNAL_19 : std_logic ;
  signal RFO2_DATA2_INTERNAL_20 : std_logic ;
  signal RFO2_DATA2_INTERNAL_21 : std_logic ;
  signal RFO2_DATA2_INTERNAL_22 : std_logic ;
  signal RFO2_DATA2_INTERNAL_23 : std_logic ;
  signal RFO2_DATA2_INTERNAL_24 : std_logic ;
  signal RFO2_DATA2_INTERNAL_25 : std_logic ;
  signal RFO2_DATA2_INTERNAL_26 : std_logic ;
  signal RFO2_DATA2_INTERNAL_27 : std_logic ;
  signal RFO2_DATA2_INTERNAL_28 : std_logic ;
  signal RFO2_DATA2_INTERNAL_29 : std_logic ;
  signal RFO2_DATA2_INTERNAL_30 : std_logic ;
  signal GND : std_logic ;
  signal VCC : std_logic ;
  signal \GRLFPC20.FPI.START\ : std_logic ;
  signal \GRLFPC20.FPI.RST_0_G0_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT\ : std_logic ;
  signal \GRLFPC20.R.I.EXEC\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY\ : std_logic ;
  signal \GRLFPC20.R.X.LD\ : std_logic ;
  signal \GRLFPC20.R.X.AFSR\ : std_logic ;
  signal \GRLFPC20.R.X.FPOP\ : std_logic ;
  signal \GRLFPC20.R.A.RS1D\ : std_logic ;
  signal \GRLFPC20.R.A.RS2D\ : std_logic ;
  signal \GRLFPC20.R.A.AFQ\ : std_logic ;
  signal \GRLFPC20.R.MK.RST\ : std_logic ;
  signal \GRLFPC20.R.MK.RST2\ : std_logic ;
  signal \GRLFPC20.R.MK.HOLDN1\ : std_logic ;
  signal \GRLFPC20.R.E.FPOP\ : std_logic ;
  signal \GRLFPC20.R.M.FPOP\ : std_logic ;
  signal \GRLFPC20.R.A.ST\ : std_logic ;
  signal \GRLFPC20.R.A.AFSR\ : std_logic ;
  signal \GRLFPC20.R.MK.HOLDN2\ : std_logic ;
  signal \GRLFPC20.R.I.V\ : std_logic ;
  signal \GRLFPC20.R.M.LD\ : std_logic ;
  signal \GRLFPC20.R.E.LD\ : std_logic ;
  signal \GRLFPC20.R.A.LD\ : std_logic ;
  signal \GRLFPC20.R.A.FPOP\ : std_logic ;
  signal \GRLFPC20.R.MK.LDOP\ : std_logic ;
  signal \GRLFPC20.R.M.AFQ\ : std_logic ;
  signal \GRLFPC20.R.M.AFSR\ : std_logic ;
  signal \GRLFPC20.R.E.AFQ\ : std_logic ;
  signal \GRLFPC20.R.E.AFSR\ : std_logic ;
  signal \GRLFPC20.R.X.AFQ\ : std_logic ;
  signal \GRLFPC20.R.A.MOV\ : std_logic ;
  signal \GRLFPC20.R.I.RDD\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY2\ : std_logic ;
  signal \GRLFPC20.R.FSR.NONSTD\ : std_logic ;
  signal \GRLFPC20.COMB.RS2D_1_IV\ : std_logic ;
  signal \GRLFPC20.COMB.V.MK.RST_1_0_G0\ : std_logic ;
  signal \GRLFPC20.RIN.MK.LDOP_X\ : std_logic ;
  signal \GRLFPC20.R.MK.HOLDN1_0_0_G0_X\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY_0_0_G0\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY2_0_0_G0_X\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_0__G0\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_2__G0\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_3__G0\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_5__G0\ : std_logic ;
  signal \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SCTRL_NEW_0_0__G0_I_M2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_4_0_2__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_5_0_1__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_0__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_65__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_18_0_74__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_374__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_375__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_114__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_0_7__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_SUM0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_26\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_47\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_20\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_26\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_45\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_38\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_61\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_58\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_61\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_19\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_58\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_59\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_60\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_61\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_19\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_59\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_61\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_19\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_46\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_52\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_53\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_15\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_41\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_46\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_58\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_61\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_24\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_24\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0_62__ROM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_45\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_56\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.CO0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_173__G0_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_172__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN38_PCTRL_NEW_I_0_G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN33_PCTRL_NEW_I_0_G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_7__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_5__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_2__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_1__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_IV_I_0_0__G0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_I_0_0__G0_0_M2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_15\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_19\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_20\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_21\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_23\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_24\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_26\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_33\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_34\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_38\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_39\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_40\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_41\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_43\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_45\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_46\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_47\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_48\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_49\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_51\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_52\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_53\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_55\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_56\ : std_logic ;
  signal N_10418 : std_logic ;
  signal N_10419 : std_logic ;
  signal N_10421 : std_logic ;
  signal N_10422 : std_logic ;
  signal N_10423 : std_logic ;
  signal N_10424 : std_logic ;
  signal N_10425 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_11\ : std_logic ;
  signal \GRLFPC20.V.STATE_0_SQMUXA_1_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G0_I_O4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_6_0_67__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_65__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_46__G2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_41__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_41__G4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_21__G2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_20__G2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_9__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_9__G4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_319__G3_0_X2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_318__G3_0_X2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_316__G3_0_X2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_258__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_112__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_112__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_111__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_111__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_110__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_110__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_109__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_109__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_108__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_108__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_107__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_107__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_106__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_106__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_105__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_105__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_104__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_104__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_103__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_103__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_102__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_102__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_101__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_101__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_100__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_100__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_99__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_99__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_98__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_98__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_97__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_97__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_96__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_96__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_95__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_95__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_94__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_94__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_93__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_93__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_92__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_92__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_91__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_91__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_90__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_90__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_89__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_89__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_88__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_88__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_87__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_87__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_86__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_86__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_85__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_85__G2_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_84__G1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_84__G2_X\ : std_logic ;
  signal \GRLFPC20.R.I.V_1_0_G3\ : std_logic ;
  signal \GRLFPC20.R.A.RDD_0_0_0__G1_0\ : std_logic ;
  signal \GRLFPC20.R.A.SEQERR_0_0_0__G1\ : std_logic ;
  signal \GRLFPC20.R.A.ST_0_0_G1\ : std_logic ;
  signal \GRLFPC20.R.A.LD_0_0_G1\ : std_logic ;
  signal \GRLFPC20.R.A.FPOP_0_0_G1\ : std_logic ;
  signal \GRLFPC20.R.A.AFSR_0_0_G1\ : std_logic ;
  signal \GRLFPC20.R.A.AFQ_0_0_G1\ : std_logic ;
  signal \GRLFPC20.COMB.RS1D_1_U\ : std_logic ;
  signal \GRLFPC20.R.FSR.NONSTD_0_0_G3_X\ : std_logic ;
  signal \GRLFPC20.R.A.MOV_0_0_G1\ : std_logic ;
  signal \GRLFPC20.R.X.LD_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.X.FPOP_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.X.AFSR_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.X.AFQ_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.M.LD_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.M.FPOP_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.M.AFSR_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.M.AFQ_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.E.LD_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.E.FPOP_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.E.AFSR_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.E.AFQ_0_0_G1_X\ : std_logic ;
  signal \GRLFPC20.R.I.CC_0_0_0__G4\ : std_logic ;
  signal \GRLFPC20.R.I.CC_0_0_1__G4\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_0__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_0__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_1__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_1__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_12__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_12__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_17__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_17__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_18__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_18__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_19__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_19__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_20__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_20__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_21__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_21__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_28__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_28__G3_X\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_29__G2\ : std_logic ;
  signal \GRLFPC20.R.E.STDATA_1_0_29__G3_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.RD_0_0_0__G3_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.RD_0_0_1__G3_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.TEM_1_0_0__G3_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.TEM_1_0_1__G3_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.TEM_1_0_2__G3_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.TEM_1_0_3__G3_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.TEM_1_0_4__G3_X\ : std_logic ;
  signal \GRLFPC20.R.STATE_0_0_0__G1\ : std_logic ;
  signal \GRLFPC20.R.STATE_0_0_1__G1\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_2__G2\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_0__G1\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_1__G1\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_2__G1\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_3__G1\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_4__G1\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_4__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.UN17_U_RDN_I_0_503_I_A2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1_520\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.UN53_SCTRL_NEW\ : std_logic ;
  signal \GRLFPC20.R.I.EXEC_0_0_G1_0_549_I\ : std_logic ;
  signal \GRLFPC20.R.I.RDD_0_0_G1_0_574_I\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_1__G2_0_624_I\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF1REN_1_670_I\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF2REN_1_734_I\ : std_logic ;
  signal RST_INTERNAL : std_logic ;
  signal \GRLFPC20.R.I.V_1_0_G0_0\ : std_logic ;
  signal \GRLFPC20.G_884\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRONEMORE\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_SUM2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.CO0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.CO0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_ANC3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.CO0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_259__G5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.COMB.WREN129\ : std_logic ;
  signal \GRLFPC20.WREN1_0_SQMUXA_1_X\ : std_logic ;
  signal \GRLFPC20.COMB.RS1_1_SN_M2_X\ : std_logic ;
  signal \GRLFPC20.R.I.V_EN_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.FSR.FCC10\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_FPCI_0_X\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_R.I.V_0\ : std_logic ;
  signal \GRLFPC20.WRADDR_0_SQMUXA_X\ : std_logic ;
  signal \GRLFPC20.WREN2_1_SQMUXA_1_1_X\ : std_logic ;
  signal \GRLFPC20.WREN2_2_SQMUXA_1\ : std_logic ;
  signal \GRLFPC20.WREN2_1_SQMUXA_1\ : std_logic ;
  signal \GRLFPC20.COMB.WREN2_11_IV\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN15_XZROUNDOUT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN23_XZROUNDOUT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN26_XZYBUSLSBS\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3\ : std_logic ;
  signal \GRLFPC20.COMB.V.STATE14\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_0__G4\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_2__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.NOTAM2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.ENTRYSHFT.S_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN6_S_0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_ENTRYPOINT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529_A3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN14_CONDITIONAL\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\ : std_logic ;
  signal \GRLFPC20.V.FSR.AEXC_2_SQMUXA\ : std_logic ;
  signal \GRLFPC20.V.FSR.AEXC_1_SQMUXA\ : std_logic ;
  signal \GRLFPC20.COMB.V.FSR.FCC10_1\ : std_logic ;
  signal \GRLFPC20.COMB.ISFPOP2_1_X\ : std_logic ;
  signal \GRLFPC20.R.STATE_0_0_0__G3\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_R.I.V\ : std_logic ;
  signal \GRLFPC20.COMB.V.STATE\ : std_logic ;
  signal \GRLFPC20.UN1_FPCI_2\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_2__G2_490\ : std_logic ;
  signal \GRLFPC20.UN1_FPCI_13\ : std_logic ;
  signal \GRLFPC20.V.STATE_1_SQMUXA_1_X\ : std_logic ;
  signal \GRLFPC20.COMB.UN7_RS1V_X\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_RS1V_X\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1.M14_0_A2_1\ : std_logic ;
  signal \GRLFPC20.R.A.RDD_0_0_0__G2\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1.M14_0_O2\ : std_logic ;
  signal \GRLFPC20.R.A.AFSR_0_0_G1_1\ : std_logic ;
  signal \GRLFPC20.COMB.QNE2\ : std_logic ;
  signal \GRLFPC20.COMB.SEQERR.UN7_OP_0_A2_X\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.LD_1_0_O2\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2\ : std_logic ;
  signal \GRLFPC20.UN1_MOV_1_SQMUXA\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.ST_0_A2\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.FPOP8_I_O3_X\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.ST3_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2_1\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.FPOP2_0_O2_X\ : std_logic ;
  signal \GRLFPC20.COMB.LOCKGEN.LOCKI_I_0_0_A2_0\ : std_logic ;
  signal \GRLFPC20.R.A.SEQERR_0_0_0__G3\ : std_logic ;
  signal \GRLFPC20.RS1D_CNST_0_A2_2_X\ : std_logic ;
  signal \GRLFPC20.COMB.RS1V_1_IV\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF1REN_1_0_650_A2_3_X\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.FPOP2_0_A2\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1.M10_2_0_A2_X\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_MEXC_1\ : std_logic ;
  signal \GRLFPC20.COMB.V.I.EXEC_5_IV\ : std_logic ;
  signal \GRLFPC20.R.I.EXC_2_0_3__G3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DECODESTATUS.UN7_STATUS\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN3_INEXACT\ : std_logic ;
  signal \GRLFPC20.COMB.ANNULRES_1_IV_454\ : std_logic ;
  signal \GRLFPC20.R.I.EXEC_0_0_G1_0_I_A8_0\ : std_logic ;
  signal \GRLFPC20.COMB.UN3_HOLDN_X\ : std_logic ;
  signal \GRLFPC20.ANNULFPU_0_SQMUXA_2_X\ : std_logic ;
  signal \GRLFPC20.COMB.V.E.STDATA2_X\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.RDD5_3_0_A2_X\ : std_logic ;
  signal \GRLFPC20.FPI.LDOP_2\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY2_0_0_G3\ : std_logic ;
  signal \GRLFPC20.ANNULRES_1_SQMUXA\ : std_logic ;
  signal \GRLFPC20.ANNULRES_0_SQMUXA_12_1\ : std_logic ;
  signal \GRLFPC20.ANNULFPU_0_SQMUXA_X\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.LD_1_0_A2_0\ : std_logic ;
  signal \GRLFPC20.COMB.RSDECODE.RS1V_X\ : std_logic ;
  signal \GRLFPC20.COMB.LOCKGEN.DEPCHECK\ : std_logic ;
  signal \GRLFPC20.ANNULFPU_0_SQMUXA_1_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_36\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTBZERODENORM\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.UN1_GRFPUS\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTAINFNAN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.UN4_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN7_SHDVAR\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8S2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTNULLEXC\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXC\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.UN2_TEMP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2_0\ : std_logic ;
  signal NN_1 : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN29_GRFPUSX_M_381\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_AREGSIGN_SEL_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT_I_M\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TEMP\ : std_logic ;
  signal \GRLFPC20.UN1_FPCI_22_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.UN17_U_RDN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.ANC1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7356\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_BNC4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_261__G5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN6_NOTPROP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.ROMXZSL2FROMC\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_STKGEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_STKOUT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN4_STKOUT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0_A3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN1_NOTPROP_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN19_GEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_2_I_O3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C1_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_43\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.RDD3_TZ\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_1_X\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.RDD4_0_A2_0_X\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.RDD4_0_A2_X\ : std_logic ;
  signal \GRLFPC20.R.A.RS1D_0_0_G4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM0\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.RDD5_0_A3\ : std_logic ;
  signal \GRLFPC20.MOV_7_SQMUXA\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF1REN_1_670_I_M4\ : std_logic ;
  signal \GRLFPC20.COMB.V.I.V_1_F1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLCREGXZ.UN1_INFORCREGDB\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_172__G0_0_M3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_AXB0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN40_SHDVAR\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0\ : std_logic ;
  signal \GRLFPC20.COMB.WREN1_11_IV\ : std_logic ;
  signal \GRLFPC20.WREN1_1_SQMUXA\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTBINFNAN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_31\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_57\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_38\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_5\ : std_logic ;
  signal \GRLFPC20.UN1_RS1V_0_SQMUXA\ : std_logic ;
  signal \GRLFPC20.RS1V_0_SQMUXA_1_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_I_O2\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_TZ\ : std_logic ;
  signal \GRLFPC20.COMB.RSDECODE.UN1_FPCI_0_X\ : std_logic ;
  signal \GRLFPC20.R.A.MOV_0_0_G1_0_X\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_0_X\ : std_logic ;
  signal \GRLFPC20.R.A.AFQ_0_0_G1_0\ : std_logic ;
  signal \GRLFPC20.V.FSR.AEXC_1_SQMUXA_0\ : std_logic ;
  signal \GRLFPC20.R.I.RDD_0_0_G1_0_574_I_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_E\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0_A2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_4\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1.M14_0_A2_0_0\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1.M14_0_A2_0_1\ : std_logic ;
  signal \GRLFPC20.R.A.AFQ_0_0_G1_0_3\ : std_logic ;
  signal \GRLFPC20.WREN1_1_SQMUXA_1\ : std_logic ;
  signal \GRLFPC20.COMB.WREN1_11_IV_1_X\ : std_logic ;
  signal \GRLFPC20.R.A.RS1D_0_0_G4_1_X\ : std_logic ;
  signal \GRLFPC20.RS2_0_SQMUXA_0_X\ : std_logic ;
  signal \GRLFPC20.UN1_MOV_1_SQMUXA_0\ : std_logic ;
  signal \GRLFPC20.COMB.LOCK_1_1_X\ : std_logic ;
  signal \GRLFPC20.MOV_2_SQMUXA_2\ : std_logic ;
  signal \GRLFPC20.RS1D_CNST_0_A2_0\ : std_logic ;
  signal \GRLFPC20.RS1D_CNST_0_A2_1_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_0__G0_0_A3_0_X\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.FPOP3_0\ : std_logic ;
  signal \GRLFPC20.COMB.RSDECODE.RS1V2_0\ : std_logic ;
  signal \GRLFPC20.COMB.WREN2_11_IV_1_X\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.UN1_FPCI_7_1_X\ : std_logic ;
  signal \GRLFPC20.R.A.MOV_0_0_G1_1_X\ : std_logic ;
  signal \GRLFPC20.R.A.MOV_0_0_G1_3\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.UN1_FPCI_0_7_2\ : std_logic ;
  signal \GRLFPC20.COMB.UN9_CCV_0_0\ : std_logic ;
  signal \GRLFPC20.COMB.UN9_CCV_0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM_0\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_A6_1_0\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_FPCI_0_1_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN4_NOTSHIFTCOUNT1_0\ : std_logic ;
  signal \GRLFPC20.N_1243_I_0_A2_1_X\ : std_logic ;
  signal \GRLFPC20.V.FSR.FTT_1_SQMUXA_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_11_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_11\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_MEXC_1_0\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_MEXC_1_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELINITREMBIT_0\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_1__G2_0_624_I_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_10\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_13\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_15\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_23\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_24\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_1_2\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN12_SRTOSTICKY_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_3_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_3\ : std_logic ;
  signal \GRLFPC20.R.A.AFSR_0_0_G1_1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN11_WQSTSETS_0\ : std_logic ;
  signal \GRLFPC20.R.STATE_0_0_0__G3_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN13_GEN_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\ : std_logic ;
  signal \GRLFPC20.R.I.EXEC_0_0_G1_0_I_0_0\ : std_logic ;
  signal \GRLFPC20.R.I.V_1_0_G0_0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_5\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_6\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_8\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_9\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_11\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_12\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_14\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_15\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_16\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_17\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_18\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_21\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_22\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_25\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_27\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_28\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_29\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_30\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_32\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_35\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_38\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_39\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_40\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_41\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_42\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_44\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_45\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_47\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_50\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_51\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_52\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_53\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_54\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M2_E_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M2_E_4\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_0__G1_0\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_3__G1_0\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_1__G1_0\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_2__G1_0\ : std_logic ;
  signal \GRLFPC20.R.FSR.AEXC_1_0_4__G1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT_I_M_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_IV_I_0_0__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_A5_0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_A5_0_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_2__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_5__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_1__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_7__G0_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_1\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY_0_0_G0_0_X\ : std_logic ;
  signal \GRLFPC20.COMB.V.MK.RST_1_0_G0_1_0_X\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\ : std_logic ;
  signal \GRLFPC20.V.FSR.CEXC_3_SQMUXA\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14S2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11S4\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_FPCI_4\ : std_logic ;
  signal \GRLFPC20.RS2_0_SQMUXA\ : std_logic ;
  signal \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\ : std_logic ;
  signal \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_R.A.RS1_1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_37\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\ : std_logic ;
  signal \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M2\ : std_logic ;
  signal \GRLFPC20.COMB.UN1_R.I.EXC\ : std_logic ;
  signal \GRLFPC20.WRADDR_1_SQMUXA\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_2\ : std_logic ;
  signal \GRLFPC20.WRADDR_0_SQMUXA_0_X\ : std_logic ;
  signal \GRLFPC20.RS1V_0_SQMUXA\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\ : std_logic ;
  signal \GRLFPC20.COMB.UN19_IUEXEC\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\ : std_logic ;
  signal \GRLFPC20.COMB.UN2_HOLDN\ : std_logic ;
  signal \GRLFPC20.V.I.EXEC_0_SQMUXA\ : std_logic ;
  signal \GRLFPC20.FPI.LDOP\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_20__G2_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M5_A\ : std_logic ;
  signal \GRLFPC20.COMB.FPDECODE.RDD3_TZ_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_0_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_1_A\ : std_logic ;
  signal \GRLFPC20.ANNULRES_1_SQMUXA_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20_A\ : std_logic ;
  signal \GRLFPC20.COMB.RDD_1.M14_0_A2_0_0_A\ : std_logic ;
  signal \GRLFPC20.COMB.RSDECODE.RS1V2_0_A\ : std_logic ;
  signal \GRLFPC20.RS1V_0_SQMUXA_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_375__G0_A\ : std_logic ;
  signal \GRLFPC20.R.MK.BUSY2_0_0_G3_A\ : std_logic ;
  signal \GRLFPC20.RS1D_CNST_0_A2_0_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_5_A\ : std_logic ;
  signal \GRLFPC20.COMB.ANNULRES_1_IV_454_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_374__G0_0_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_9_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_35_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_114__G0_A\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_S\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_6_0_67__G0_E_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\ : std_logic ;
  signal \GRLFPC20.R.I.PC_1_0_2__G2_X_I\ : std_logic ;
  signal \GRLFPC20.R.FSR.FTT_1_0_0__G0_I_O4_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2_RETI\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_RETI\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1_RETI\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES_RETI\ : std_logic ;
  signal N_19146 : std_logic ;
  signal N_19147 : std_logic ;
  signal N_19148 : std_logic ;
  signal N_19149 : std_logic ;
  signal N_19200 : std_logic ;
  signal N_19201 : std_logic ;
  signal N_19202 : std_logic ;
  signal N_19203 : std_logic ;
  signal N_19204 : std_logic ;
  signal N_19205 : std_logic ;
  signal N_19206 : std_logic ;
  signal N_19207 : std_logic ;
  signal N_19208 : std_logic ;
  signal N_19209 : std_logic ;
  signal N_19210 : std_logic ;
  signal N_19211 : std_logic ;
  signal N_19212 : std_logic ;
  signal N_19213 : std_logic ;
  signal N_19214 : std_logic ;
  signal N_19215 : std_logic ;
  signal N_19216 : std_logic ;
  signal N_19217 : std_logic ;
  signal N_19218 : std_logic ;
  signal N_19219 : std_logic ;
  signal N_19220 : std_logic ;
  signal N_19221 : std_logic ;
  signal N_19222 : std_logic ;
  signal N_19223 : std_logic ;
  signal N_19224 : std_logic ;
  signal N_19225 : std_logic ;
  signal N_19226 : std_logic ;
  signal N_19227 : std_logic ;
  signal N_19228 : std_logic ;
  signal N_19229 : std_logic ;
  signal N_19230 : std_logic ;
  signal N_19231 : std_logic ;
  signal N_19232 : std_logic ;
  signal N_19233 : std_logic ;
  signal N_19234 : std_logic ;
  signal N_19235 : std_logic ;
  signal N_19236 : std_logic ;
  signal N_19237 : std_logic ;
  signal N_19238 : std_logic ;
  signal N_19239 : std_logic ;
  signal N_19240 : std_logic ;
  signal N_19241 : std_logic ;
  signal N_19242 : std_logic ;
  signal N_19243 : std_logic ;
  signal N_19244 : std_logic ;
  signal N_19245 : std_logic ;
  signal N_19246 : std_logic ;
  signal N_19247 : std_logic ;
  signal N_19248 : std_logic ;
  signal N_19249 : std_logic ;
  signal N_19250 : std_logic ;
  signal N_19251 : std_logic ;
  signal N_19252 : std_logic ;
  signal N_19253 : std_logic ;
  signal N_19254 : std_logic ;
  signal N_19255 : std_logic ;
  signal N_19256 : std_logic ;
  signal N_19257 : std_logic ;
  signal N_19258 : std_logic ;
  signal N_19259 : std_logic ;
  signal N_19260 : std_logic ;
  signal N_19261 : std_logic ;
  signal N_19262 : std_logic ;
  signal N_19263 : std_logic ;
  signal N_19264 : std_logic ;
  signal N_19265 : std_logic ;
  signal N_19266 : std_logic ;
  signal N_19267 : std_logic ;
  signal N_19268 : std_logic ;
  signal N_19269 : std_logic ;
  signal N_19270 : std_logic ;
  signal N_19271 : std_logic ;
  signal N_19272 : std_logic ;
  signal N_19273 : std_logic ;
  signal N_19274 : std_logic ;
  signal N_19275 : std_logic ;
  signal N_19276 : std_logic ;
  signal N_19277 : std_logic ;
  signal N_19278 : std_logic ;
  signal N_19279 : std_logic ;
  signal N_19280 : std_logic ;
  signal N_19281 : std_logic ;
  signal N_19282 : std_logic ;
  signal N_19283 : std_logic ;
  signal N_19284 : std_logic ;
  signal N_19285 : std_logic ;
  signal N_19286 : std_logic ;
  signal N_19287 : std_logic ;
  signal N_19288 : std_logic ;
  signal N_19289 : std_logic ;
  signal N_19290 : std_logic ;
  signal N_19291 : std_logic ;
  signal N_19292 : std_logic ;
  signal N_19293 : std_logic ;
  signal N_19294 : std_logic ;
  signal N_19295 : std_logic ;
  signal N_19296 : std_logic ;
  signal N_19297 : std_logic ;
  signal N_19298 : std_logic ;
  signal N_19299 : std_logic ;
  signal N_19300 : std_logic ;
  signal N_19301 : std_logic ;
  signal N_19302 : std_logic ;
  signal N_19303 : std_logic ;
  signal N_19304 : std_logic ;
  signal N_19305 : std_logic ;
  signal N_19306 : std_logic ;
  signal N_27907 : std_logic ;
  signal N_27908 : std_logic ;
  signal HOLDN_INTERNAL : std_logic ;
  signal CPI_DBG_FSR_INTERNAL : std_logic ;
  signal CPI_DBG_ADDR_INTERNAL : std_logic ;
  signal N_1 : std_logic ;
  signal N_2 : std_logic ;
  signal N_3 : std_logic ;
  signal N_4 : std_logic ;
  signal N_5 : std_logic ;
  signal N_6 : std_logic ;
  signal N_7 : std_logic ;
  signal N_8 : std_logic ;
  signal N_9 : std_logic ;
  signal N_10 : std_logic ;
  signal N_11 : std_logic ;
  signal N_12 : std_logic ;
  signal N_13 : std_logic ;
  signal N_14 : std_logic ;
  signal N_15 : std_logic ;
  signal N_16 : std_logic ;
  signal N_17 : std_logic ;
  signal N_18 : std_logic ;
  signal N_19 : std_logic ;
  signal N_20 : std_logic ;
  signal N_21 : std_logic ;
  signal N_22 : std_logic ;
  signal N_23 : std_logic ;
  signal N_24 : std_logic ;
  signal N_25 : std_logic ;
  signal N_26 : std_logic ;
  signal N_27 : std_logic ;
  signal N_28 : std_logic ;
  signal N_29 : std_logic ;
  signal N_30 : std_logic ;
  signal N_31 : std_logic ;
  signal N_32 : std_logic ;
  signal N_33 : std_logic ;
  signal N_34 : std_logic ;
  signal N_35 : std_logic ;
  signal N_36 : std_logic ;
  signal N_37 : std_logic ;
  signal N_38 : std_logic ;
  signal N_39 : std_logic ;
  signal N_40 : std_logic ;
  signal N_41 : std_logic ;
  signal N_42 : std_logic ;
  signal N_43 : std_logic ;
  signal N_44 : std_logic ;
  signal N_45 : std_logic ;
  signal N_46 : std_logic ;
  signal N_47 : std_logic ;
  signal N_48 : std_logic ;
  signal N_49 : std_logic ;
  signal N_50 : std_logic ;
  signal N_51 : std_logic ;
  signal N_52 : std_logic ;
  signal N_53 : std_logic ;
  signal N_54 : std_logic ;
  signal N_55 : std_logic ;
  signal N_56 : std_logic ;
  signal N_57 : std_logic ;
  signal N_58 : std_logic ;
  signal N_59 : std_logic ;
  signal N_60 : std_logic ;
  signal N_61 : std_logic ;
  signal N_62 : std_logic ;
  signal N_63 : std_logic ;
  signal N_64 : std_logic ;
  signal N_65 : std_logic ;
  signal N_66 : std_logic ;
  signal N_67 : std_logic ;
  signal N_68 : std_logic ;
  signal N_69 : std_logic ;
  signal N_70 : std_logic ;
  signal N_71 : std_logic ;
  signal N_72 : std_logic ;
  signal N_73 : std_logic ;
  signal N_74 : std_logic ;
  signal N_75 : std_logic ;
  signal N_76 : std_logic ;
  signal N_77 : std_logic ;
  signal N_78 : std_logic ;
  signal N_79 : std_logic ;
  signal N_80 : std_logic ;
  signal N_81 : std_logic ;
  signal N_82 : std_logic ;
  signal N_83 : std_logic ;
  signal N_84 : std_logic ;
  signal N_85 : std_logic ;
  signal N_86 : std_logic ;
  signal N_87 : std_logic ;
  signal N_88 : std_logic ;
  signal N_89 : std_logic ;
  signal N_90 : std_logic ;
  signal N_91 : std_logic ;
  signal N_92 : std_logic ;
  signal N_93 : std_logic ;
  signal N_94 : std_logic ;
  signal N_95 : std_logic ;
  signal N_96 : std_logic ;
  signal N_97 : std_logic ;
  signal N_98 : std_logic ;
  signal N_99 : std_logic ;
  signal N_100 : std_logic ;
  signal N_101 : std_logic ;
  signal N_102 : std_logic ;
  signal N_103 : std_logic ;
  signal N_104 : std_logic ;
  signal N_105 : std_logic ;
  signal N_106 : std_logic ;
  signal N_107 : std_logic ;
  signal N_108 : std_logic ;
  signal N_109 : std_logic ;
  signal N_110 : std_logic ;
  signal N_111 : std_logic ;
  signal N_112 : std_logic ;
  signal N_113 : std_logic ;
  signal N_114 : std_logic ;
  signal N_115 : std_logic ;
  signal N_116 : std_logic ;
  signal N_117 : std_logic ;
  signal N_118 : std_logic ;
  signal N_119 : std_logic ;
  signal N_120 : std_logic ;
  signal N_121 : std_logic ;
  signal N_122 : std_logic ;
  signal N_123 : std_logic ;
  signal N_124 : std_logic ;
  signal N_125 : std_logic ;
  signal N_126 : std_logic ;
  signal N_127 : std_logic ;
  signal N_128 : std_logic ;
  signal N_129 : std_logic ;
  signal N_130 : std_logic ;
  signal N_131 : std_logic ;
  signal N_132 : std_logic ;
  signal N_133 : std_logic ;
  signal N_134 : std_logic ;
  signal N_135 : std_logic ;
  signal N_136 : std_logic ;
  signal N_137 : std_logic ;
  signal N_138 : std_logic ;
  signal N_139 : std_logic ;
  signal N_140 : std_logic ;
  signal N_141 : std_logic ;
  signal N_142 : std_logic ;
  signal N_143 : std_logic ;
  signal N_144 : std_logic ;
  signal N_145 : std_logic ;
  signal N_146 : std_logic ;
  signal N_147 : std_logic ;
  signal N_148 : std_logic ;
  signal N_149 : std_logic ;
  signal N_150 : std_logic ;
  signal N_151 : std_logic ;
  signal N_152 : std_logic ;
  signal N_153 : std_logic ;
  signal N_154 : std_logic ;
  signal N_155 : std_logic ;
  signal N_156 : std_logic ;
  signal N_157 : std_logic ;
  signal N_158 : std_logic ;
  signal N_159 : std_logic ;
  signal N_160 : std_logic ;
  signal N_161 : std_logic ;
  signal N_162 : std_logic ;
  signal N_163 : std_logic ;
  signal N_164 : std_logic ;
  signal N_165 : std_logic ;
  signal N_166 : std_logic ;
  signal N_167 : std_logic ;
  signal N_168 : std_logic ;
  signal N_169 : std_logic ;
  signal N_170 : std_logic ;
  signal N_171 : std_logic ;
  signal N_172 : std_logic ;
  signal N_173 : std_logic ;
  signal N_174 : std_logic ;
  signal N_175 : std_logic ;
  signal N_176 : std_logic ;
  signal N_177 : std_logic ;
  signal N_178 : std_logic ;
  signal N_179 : std_logic ;
  signal N_180 : std_logic ;
  signal N_181 : std_logic ;
  signal N_182 : std_logic ;
  signal N_183 : std_logic ;
  signal N_184 : std_logic ;
  signal N_185 : std_logic ;
  signal N_186 : std_logic ;
  signal N_187 : std_logic ;
  signal N_188 : std_logic ;
  signal N_189 : std_logic ;
  signal N_190 : std_logic ;
  signal N_191 : std_logic ;
  signal N_192 : std_logic ;
  signal N_193 : std_logic ;
  signal N_194 : std_logic ;
  signal N_195 : std_logic ;
  signal N_196 : std_logic ;
  signal N_197 : std_logic ;
  signal N_198 : std_logic ;
  signal N_199 : std_logic ;
  signal N_200 : std_logic ;
  signal N_201 : std_logic ;
  signal N_202 : std_logic ;
  signal N_203 : std_logic ;
  signal N_204 : std_logic ;
  signal N_205 : std_logic ;
  signal N_206 : std_logic ;
  signal N_207 : std_logic ;
  signal N_208 : std_logic ;
  signal N_209 : std_logic ;
  signal N_210 : std_logic ;
  signal N_211 : std_logic ;
  signal N_212 : std_logic ;
  signal N_213 : std_logic ;
  signal N_214 : std_logic ;
  signal N_215 : std_logic ;
  signal N_216 : std_logic ;
  signal N_217 : std_logic ;
  signal N_218 : std_logic ;
  signal N_219 : std_logic ;
  signal N_220 : std_logic ;
  signal N_221 : std_logic ;
  signal N_222 : std_logic ;
  signal N_223 : std_logic ;
  signal N_224 : std_logic ;
  signal N_225 : std_logic ;
  signal N_226 : std_logic ;
  signal N_227 : std_logic ;
  signal N_228 : std_logic ;
  signal N_229 : std_logic ;
  signal N_230 : std_logic ;
  signal N_231 : std_logic ;
  signal N_232 : std_logic ;
  signal N_233 : std_logic ;
  signal N_234 : std_logic ;
  signal N_235 : std_logic ;
  signal N_236 : std_logic ;
  signal N_237 : std_logic ;
  signal N_238 : std_logic ;
  signal N_239 : std_logic ;
  signal N_240 : std_logic ;
  signal N_241 : std_logic ;
  signal N_242 : std_logic ;
  signal N_243 : std_logic ;
  signal N_244 : std_logic ;
  signal N_245 : std_logic ;
  signal N_246 : std_logic ;
  signal N_247 : std_logic ;
  signal N_248 : std_logic ;
  signal N_249 : std_logic ;
  signal N_250 : std_logic ;
  signal N_251 : std_logic ;
  signal N_252 : std_logic ;
  signal N_253 : std_logic ;
  signal N_254 : std_logic ;
  signal N_255 : std_logic ;
  signal N_256 : std_logic ;
  signal N_257 : std_logic ;
  signal N_258 : std_logic ;
  signal N_259 : std_logic ;
  signal N_260 : std_logic ;
  signal N_261 : std_logic ;
  signal N_262 : std_logic ;
  signal N_263 : std_logic ;
  signal N_264 : std_logic ;
  signal N_265 : std_logic ;
  signal N_266 : std_logic ;
  signal N_267 : std_logic ;
  signal N_268 : std_logic ;
  signal N_269 : std_logic ;
  signal N_270 : std_logic ;
  signal N_271 : std_logic ;
  signal N_272 : std_logic ;
  signal N_273 : std_logic ;
  signal N_274 : std_logic ;
  signal N_275 : std_logic ;
  signal N_276 : std_logic ;
  signal N_277 : std_logic ;
  signal N_278 : std_logic ;
  signal N_279 : std_logic ;
  signal N_280 : std_logic ;
  signal N_281 : std_logic ;
  signal N_282 : std_logic ;
  signal N_283 : std_logic ;
  signal N_284 : std_logic ;
  signal N_285 : std_logic ;
  signal N_286 : std_logic ;
  signal N_287 : std_logic ;
  signal N_288 : std_logic ;
  signal N_289 : std_logic ;
  signal N_290 : std_logic ;
  signal N_291 : std_logic ;
  signal N_292 : std_logic ;
  signal N_293 : std_logic ;
  signal N_294 : std_logic ;
  signal N_295 : std_logic ;
  signal N_296 : std_logic ;
  signal N_297 : std_logic ;
  signal N_298 : std_logic ;
  signal N_299 : std_logic ;
  signal N_300 : std_logic ;
  signal N_301 : std_logic ;
  signal N_302 : std_logic ;
  signal N_303 : std_logic ;
  signal N_304 : std_logic ;
  signal N_305 : std_logic ;
  signal N_306 : std_logic ;
  signal N_307 : std_logic ;
  signal N_308 : std_logic ;
  signal N_309 : std_logic ;
  signal N_310 : std_logic ;
  signal N_311 : std_logic ;
  signal N_312 : std_logic ;
  signal N_313 : std_logic ;
  signal N_314 : std_logic ;
  signal N_315 : std_logic ;
  signal N_316 : std_logic ;
  signal N_317 : std_logic ;
  signal N_318 : std_logic ;
  signal N_319 : std_logic ;
  signal N_320 : std_logic ;
  signal N_321 : std_logic ;
  signal N_322 : std_logic ;
  signal N_323 : std_logic ;
  signal N_324 : std_logic ;
  signal N_325 : std_logic ;
  signal N_326 : std_logic ;
  signal N_327 : std_logic ;
  signal N_328 : std_logic ;
  signal N_329 : std_logic ;
  signal N_330 : std_logic ;
  signal N_331 : std_logic ;
  signal N_332 : std_logic ;
  signal N_333 : std_logic ;
  signal N_334 : std_logic ;
  signal N_335 : std_logic ;
  signal N_336 : std_logic ;
  signal N_337 : std_logic ;
  signal N_338 : std_logic ;
  signal N_339 : std_logic ;
  signal N_340 : std_logic ;
  signal N_341 : std_logic ;
  signal N_342 : std_logic ;
  signal N_343 : std_logic ;
  signal N_344 : std_logic ;
  signal N_345 : std_logic ;
  signal N_346 : std_logic ;
  signal N_347 : std_logic ;
  signal N_348 : std_logic ;
  signal N_349 : std_logic ;
  signal N_350 : std_logic ;
  signal N_351 : std_logic ;
  signal N_352 : std_logic ;
  signal N_353 : std_logic ;
  signal N_354 : std_logic ;
  signal N_355 : std_logic ;
  signal N_356 : std_logic ;
  signal N_357 : std_logic ;
  signal N_358 : std_logic ;
  signal N_359 : std_logic ;
  signal N_360 : std_logic ;
  signal N_361 : std_logic ;
  signal N_362 : std_logic ;
  signal N_363 : std_logic ;
  signal N_364 : std_logic ;
  signal N_365 : std_logic ;
  signal N_366 : std_logic ;
  signal N_367 : std_logic ;
  signal N_368 : std_logic ;
  signal N_369 : std_logic ;
  signal N_370 : std_logic ;
  signal N_371 : std_logic ;
  signal N_372 : std_logic ;
  signal N_373 : std_logic ;
  signal N_374 : std_logic ;
  signal N_375 : std_logic ;
  signal N_376 : std_logic ;
  signal N_377 : std_logic ;
  signal N_378 : std_logic ;
  signal N_379 : std_logic ;
  signal N_380 : std_logic ;
  signal N_381 : std_logic ;
  signal N_382 : std_logic ;
  signal N_383 : std_logic ;
  signal N_384 : std_logic ;
  signal N_385 : std_logic ;
  signal N_386 : std_logic ;
  signal N_387 : std_logic ;
  signal N_388 : std_logic ;
  signal N_389 : std_logic ;
  signal N_390 : std_logic ;
  signal N_391 : std_logic ;
  signal N_392 : std_logic ;
  signal N_393 : std_logic ;
  signal N_394 : std_logic ;
  signal N_395 : std_logic ;
  signal N_396 : std_logic ;
  signal N_397 : std_logic ;
  signal N_398 : std_logic ;
  signal N_399 : std_logic ;
  signal N_400 : std_logic ;
  signal N_401 : std_logic ;
  signal N_402 : std_logic ;
  signal N_403 : std_logic ;
  signal N_404 : std_logic ;
  signal N_405 : std_logic ;
  signal N_406 : std_logic ;
  signal N_407 : std_logic ;
  signal N_408 : std_logic ;
  signal N_409 : std_logic ;
  signal N_410 : std_logic ;
  signal N_411 : std_logic ;
  signal N_412 : std_logic ;
  signal N_413 : std_logic ;
  signal N_414 : std_logic ;
  signal N_415 : std_logic ;
  signal N_416 : std_logic ;
  signal N_417 : std_logic ;
  signal N_418 : std_logic ;
  signal N_419 : std_logic ;
  signal N_420 : std_logic ;
  signal N_421 : std_logic ;
  signal N_422 : std_logic ;
  signal N_423 : std_logic ;
  signal N_424 : std_logic ;
  signal N_425 : std_logic ;
  signal N_426 : std_logic ;
  signal N_427 : std_logic ;
  signal N_0 : std_logic ;
  signal N_1_0 : std_logic ;
  signal N_2_0 : std_logic ;
  signal N_3_0 : std_logic ;
  signal N_4_0 : std_logic ;
  signal N_5_0 : std_logic ;
  signal N_6_0 : std_logic ;
  signal N_7_0 : std_logic ;
  signal N_8_0 : std_logic ;
  signal N_9_0 : std_logic ;
  signal N_10_0 : std_logic ;
  signal N_11_0 : std_logic ;
  signal N_12_0 : std_logic ;
  signal N_13_0 : std_logic ;
  signal N_14_0 : std_logic ;
  signal N_15_0 : std_logic ;
  signal N_16_0 : std_logic ;
  signal N_17_0 : std_logic ;
  signal N_18_0 : std_logic ;
  signal N_19_0 : std_logic ;
  signal N_20_0 : std_logic ;
  signal N_21_0 : std_logic ;
  signal N_22_0 : std_logic ;
  signal N_23_0 : std_logic ;
  signal N_24_0 : std_logic ;
  signal N_25_0 : std_logic ;
  signal N_26_0 : std_logic ;
  signal N_27_0 : std_logic ;
  signal N_28_0 : std_logic ;
  signal N_29_0 : std_logic ;
  signal N_30_0 : std_logic ;
  signal N_31_0 : std_logic ;
  signal N_32_0 : std_logic ;
  signal N_33_0 : std_logic ;
  signal N_34_0 : std_logic ;
  signal N_35_0 : std_logic ;
  signal N_36_0 : std_logic ;
  signal N_37_0 : std_logic ;
  signal N_38_0 : std_logic ;
  signal N_39_0 : std_logic ;
  signal N_40_0 : std_logic ;
  signal N_41_0 : std_logic ;
  signal N_42_0 : std_logic ;
  signal N_43_0 : std_logic ;
  signal N_44_0 : std_logic ;
  signal N_45_0 : std_logic ;
  signal N_46_0 : std_logic ;
  signal N_47_0 : std_logic ;
  signal N_48_0 : std_logic ;
  signal N_49_0 : std_logic ;
  signal N_50_0 : std_logic ;
  signal N_51_0 : std_logic ;
  signal N_52_0 : std_logic ;
  signal N_53_0 : std_logic ;
  signal N_54_0 : std_logic ;
  signal N_55_0 : std_logic ;
  signal N_56_0 : std_logic ;
  signal N_57_0 : std_logic ;
  signal N_58_0 : std_logic ;
  signal N_59_0 : std_logic ;
  signal N_60_0 : std_logic ;
  signal N_61_0 : std_logic ;
  signal N_62_0 : std_logic ;
  signal N_63_0 : std_logic ;
  signal N_64_0 : std_logic ;
  signal N_65_0 : std_logic ;
  signal N_66_0 : std_logic ;
  signal N_67_0 : std_logic ;
  signal N_68_0 : std_logic ;
  signal N_69_0 : std_logic ;
  signal N_70_0 : std_logic ;
  signal N_71_0 : std_logic ;
  signal N_72_0 : std_logic ;
  signal N_73_0 : std_logic ;
  signal N_74_0 : std_logic ;
  signal N_75_0 : std_logic ;
  signal N_76_0 : std_logic ;
  signal N_77_0 : std_logic ;
  signal N_78_0 : std_logic ;
  signal N_79_0 : std_logic ;
  signal N_80_0 : std_logic ;
  signal N_81_0 : std_logic ;
  signal N_82_0 : std_logic ;
  signal N_83_0 : std_logic ;
  signal N_84_0 : std_logic ;
  signal N_85_0 : std_logic ;
  signal N_86_0 : std_logic ;
  signal N_87_0 : std_logic ;
  signal N_88_0 : std_logic ;
  signal N_89_0 : std_logic ;
  signal N_90_0 : std_logic ;
  signal N_91_0 : std_logic ;
  signal N_92_0 : std_logic ;
  signal N_93_0 : std_logic ;
  signal N_94_0 : std_logic ;
  signal N_95_0 : std_logic ;
  signal N_96_0 : std_logic ;
  signal N_97_0 : std_logic ;
  signal N_98_0 : std_logic ;
  signal N_99_0 : std_logic ;
  signal N_100_0 : std_logic ;
  signal N_101_0 : std_logic ;
  signal N_102_0 : std_logic ;
  signal N_103_0 : std_logic ;
  signal N_104_0 : std_logic ;
  signal N_105_0 : std_logic ;
  signal N_106_0 : std_logic ;
  signal N_107_0 : std_logic ;
  signal N_108_0 : std_logic ;
  signal N_109_0 : std_logic ;
  signal N_110_0 : std_logic ;
  signal N_111_0 : std_logic ;
  signal N_112_0 : std_logic ;
  signal N_113_0 : std_logic ;
  signal N_114_0 : std_logic ;
  signal N_115_0 : std_logic ;
  signal N_116_0 : std_logic ;
  signal N_117_0 : std_logic ;
  signal N_118_0 : std_logic ;
  signal N_119_0 : std_logic ;
  signal N_120_0 : std_logic ;
  signal N_121_0 : std_logic ;
  signal N_122_0 : std_logic ;
  signal N_123_0 : std_logic ;
  signal N_124_0 : std_logic ;
  signal N_125_0 : std_logic ;
  signal N_126_0 : std_logic ;
  signal N_127_0 : std_logic ;
  signal N_128_0 : std_logic ;
  signal N_129_0 : std_logic ;
  signal N_130_0 : std_logic ;
  signal N_131_0 : std_logic ;
  signal N_132_0 : std_logic ;
  signal N_133_0 : std_logic ;
  signal N_134_0 : std_logic ;
  signal N_135_0 : std_logic ;
  signal N_136_0 : std_logic ;
  signal N_137_0 : std_logic ;
  signal N_138_0 : std_logic ;
  signal N_139_0 : std_logic ;
  signal N_140_0 : std_logic ;
  signal N_141_0 : std_logic ;
  signal N_142_0 : std_logic ;
  signal N_143_0 : std_logic ;
  signal N_144_0 : std_logic ;
  signal N_145_0 : std_logic ;
  signal N_146_0 : std_logic ;
  signal N_147_0 : std_logic ;
  signal N_148_0 : std_logic ;
  signal N_149_0 : std_logic ;
  signal N_150_0 : std_logic ;
  signal N_151_0 : std_logic ;
  signal N_152_0 : std_logic ;
  signal N_153_0 : std_logic ;
  signal N_154_0 : std_logic ;
  signal N_155_0 : std_logic ;
  signal N_156_0 : std_logic ;
  signal N_157_0 : std_logic ;
  signal N_158_0 : std_logic ;
  signal N_159_0 : std_logic ;
  signal N_160_0 : std_logic ;
  signal N_161_0 : std_logic ;
  signal N_162_0 : std_logic ;
  signal N_163_0 : std_logic ;
  signal N_592 : std_logic ;
  signal N_593 : std_logic ;
  signal N_594 : std_logic ;
  signal N_595 : std_logic ;
  signal N_596 : std_logic ;
  signal N_597 : std_logic ;
  signal N_598 : std_logic ;
  signal N_599 : std_logic ;
  signal N_600 : std_logic ;
  signal N_601 : std_logic ;
  signal N_602 : std_logic ;
  signal N_603 : std_logic ;
  signal N_604 : std_logic ;
  signal N_605 : std_logic ;
  signal N_606 : std_logic ;
  signal N_607 : std_logic ;
  signal N_608 : std_logic ;
  signal N_609 : std_logic ;
  signal N_610 : std_logic ;
  signal N_611 : std_logic ;
  signal N_612 : std_logic ;
  signal N_613 : std_logic ;
  signal N_614 : std_logic ;
  signal N_615 : std_logic ;
  signal N_616 : std_logic ;
  signal N_617 : std_logic ;
  signal N_618 : std_logic ;
  signal N_619 : std_logic ;
  signal N_620 : std_logic ;
  signal N_621 : std_logic ;
  signal N_622 : std_logic ;
  signal N_623 : std_logic ;
  signal N_624 : std_logic ;
  signal N_625 : std_logic ;
  signal N_626 : std_logic ;
  signal N_627 : std_logic ;
  signal N_628 : std_logic ;
  signal N_629 : std_logic ;
  signal N_630 : std_logic ;
  signal N_631 : std_logic ;
  signal N_632 : std_logic ;
  signal N_633 : std_logic ;
  signal N_634 : std_logic ;
  signal N_635 : std_logic ;
  signal N_636 : std_logic ;
  signal N_637 : std_logic ;
  signal N_638 : std_logic ;
  signal N_639 : std_logic ;
  signal N_640 : std_logic ;
  signal N_641 : std_logic ;
  signal N_642 : std_logic ;
  signal N_643 : std_logic ;
  signal N_644 : std_logic ;
  signal N_645 : std_logic ;
  signal N_646 : std_logic ;
  signal N_647 : std_logic ;
  signal N_648 : std_logic ;
  signal N_649 : std_logic ;
  signal N_650 : std_logic ;
  signal N_651 : std_logic ;
  signal N_652 : std_logic ;
  signal N_653 : std_logic ;
  signal N_654 : std_logic ;
  signal N_655 : std_logic ;
  signal N_656 : std_logic ;
  signal N_657 : std_logic ;
  signal N_658 : std_logic ;
  signal N_659 : std_logic ;
  signal N_660 : std_logic ;
  signal N_661 : std_logic ;
  signal N_662 : std_logic ;
  signal N_663 : std_logic ;
  signal N_664 : std_logic ;
  signal N_665 : std_logic ;
  signal N_666 : std_logic ;
  signal N_667 : std_logic ;
  signal N_668 : std_logic ;
  signal N_669 : std_logic ;
  signal N_670 : std_logic ;
  signal N_671 : std_logic ;
  signal N_672 : std_logic ;
  signal N_673 : std_logic ;
  signal N_674 : std_logic ;
  signal N_675 : std_logic ;
  signal N_676 : std_logic ;
  signal N_677 : std_logic ;
  signal N_678 : std_logic ;
  signal N_679 : std_logic ;
  signal N_680 : std_logic ;
  signal N_681 : std_logic ;
  signal N_682 : std_logic ;
  signal N_683 : std_logic ;
  signal N_684 : std_logic ;
  signal N_685 : std_logic ;
  signal N_686 : std_logic ;
  signal N_687 : std_logic ;
  signal N_688 : std_logic ;
  signal N_689 : std_logic ;
  signal N_690 : std_logic ;
  signal N_691 : std_logic ;
  signal N_692 : std_logic ;
  signal N_693 : std_logic ;
  signal N_694 : std_logic ;
  signal N_695 : std_logic ;
  signal N_696 : std_logic ;
  signal N_697 : std_logic ;
  signal N_698 : std_logic ;
  signal N_699 : std_logic ;
  signal N_700 : std_logic ;
  signal N_701 : std_logic ;
  signal N_702 : std_logic ;
  signal N_703 : std_logic ;
  signal N_704 : std_logic ;
  signal N_705 : std_logic ;
  signal N_706 : std_logic ;
  signal N_707 : std_logic ;
  signal N_708 : std_logic ;
  signal N_709 : std_logic ;
  signal N_710 : std_logic ;
  signal N_711 : std_logic ;
  signal N_712 : std_logic ;
  signal N_713 : std_logic ;
  signal N_714 : std_logic ;
  signal N_715 : std_logic ;
  signal N_716 : std_logic ;
  signal N_717 : std_logic ;
  signal N_718 : std_logic ;
  signal N_719 : std_logic ;
  signal N_1_I : std_logic ;
  signal \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\ : std_logic ;
  signal \GRLFPC20.V.I.EXEC_0_SQMUXA_I\ : std_logic ;
  signal \GRLFPC20.R.A.AFQ_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\ : std_logic ;
  signal \GRLFPC20.FPI.LDOP_I\ : std_logic ;
  signal \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\ : std_logic ;
  signal \GRLFPC20.COMB.UN2_HOLDN_I\ : std_logic ;
  signal CPO_EXCZ : std_logic ;
  signal CPO_CCVZ : std_logic ;
  signal CPO_LDLOCKZ : std_logic ;
  signal CPO_HOLDNZ : std_logic ;
  signal RFI1_REN1Z : std_logic ;
  signal RFI1_REN2Z : std_logic ;
  signal RFI1_WRENZ : std_logic ;
  signal RFI2_REN1Z : std_logic ;
  signal RFI2_REN2Z : std_logic ;
  signal RFI2_WRENZ : std_logic ;
begin
GND <= '0';
VCC <= '1';
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNID87_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19306,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(20));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_RNIMEBFA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(98),
cin => N_19305);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNILF6_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19304,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(19));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1_RNIN1F1A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(99),
cin => N_19303);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIKE6_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19302,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(18));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_RNIF46C9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(100),
cin => N_19301);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIJD6_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19300,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(17));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_RNI4J5P8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(101),
cin => N_19299);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIIC6_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19298,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(16));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_RNINUSR8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(102),
cin => N_19297);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHB6_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19296,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(15));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_RNIV9EK8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(103),
cin => N_19295);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGA6_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19294,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(14));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1_RNIB5F09_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(104),
cin => N_19293);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIF96_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19292,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(13));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_RNIMGO99_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(105),
cin => N_19291);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIE86_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19290,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(12));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1_RNI6C739_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(106),
cin => N_19289);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNID76_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19288,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(11));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2_RNIR4PF8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(107),
cin => N_19287);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIC66_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19286,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(10));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_RNIIBQE8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(108),
cin => N_19285);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI4UHE_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19284,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(9));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_RNIBESB8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(109),
cin => N_19283);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI3THE_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19282,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(8));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_RNIV6LT8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(110),
cin => N_19281);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI2SHE_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19280,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(7));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3_RNIS0B5A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(111),
cin => N_19279);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNI1RHE_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19278,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(6));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2_RNIHPCSA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(112),
cin => N_19277);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIJF8_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19276,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(35));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_RNI19488_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(83),
cin => N_19275);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIIE8_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19274,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(34));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_RNIUDDV8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(84),
cin => N_19273);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHD8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19272,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(33));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_RNIED6P8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(85),
cin => N_19271);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGC8_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19270,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(32));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_RNIBDC59_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(86),
cin => N_19269);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIFB8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19268,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(31));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_RNIK7719_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(87),
cin => N_19267);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIEA8_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19266,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(30));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2_RNITT8G9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(88),
cin => N_19265);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIMH7_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19264,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(29));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1_RNIIIT0A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(89),
cin => N_19263);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNILG7_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19262,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(28));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_RNISAPE9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(90),
cin => N_19261);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIKF7_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19260,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(27));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3_RNI7TJD9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(91),
cin => N_19259);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIJE7_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19258,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(26));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_RNIKVCQ9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(92),
cin => N_19257);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIID7_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19256,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(25));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1_RNIV0RCA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(93),
cin => N_19255);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHC7_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19254,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(24));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1_RNIDGMNA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(94),
cin => N_19253);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGB7_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19252,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(23));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_RNI0404A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(95),
cin => N_19251);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIFA7_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19250,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(22));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_RNIS09P9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(96),
cin => N_19249);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIE97_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19248,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(21));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2_RNIS4ES9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(97),
cin => N_19247);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGEA_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19246,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(50));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2_RNI1SQT8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(68),
cin => N_19245);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIOL9_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19244,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(49));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3_RNIVTLE9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(69),
cin => N_19243);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNINK9_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19242,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(48));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3_RNIC4DV9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(70),
cin => N_19241);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIMJ9_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19240,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(47));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_RNIPU129_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(71),
cin => N_19239);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNILI9_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19238,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(46));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_RNITQ8H8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(72),
cin => N_19237);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIKH9_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19236,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(45));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_RNI2QIA8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(73),
cin => N_19235);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIJG9_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19234,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(44));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1_RNI4MR69_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(74),
cin => N_19233);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIIF9_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19232,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(43));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2_RNIMAHU9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(75),
cin => N_19231);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHE9_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19230,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(42));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3_RNI4RA0A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(76),
cin => N_19229);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIGD9_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19228,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(41));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1_RNIOGM2A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(77),
cin => N_19227);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIFC9_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19226,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(40));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_RNIOP1MA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(78),
cin => N_19225);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNINJ8_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19224,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(39));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_RNI5SV2A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(79),
cin => N_19223);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIMI8_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19222,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(38));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3_RNIV0AK9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(80),
cin => N_19221);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNILH8_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19220,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(37));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_RNI86OH8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(81),
cin => N_19219);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIKG8_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19218,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(36));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2_RNI90IR7_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(82),
cin => N_19217);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNINLA_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19216,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_RNIMIFAC_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(61),
cin => N_19215);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIMKA_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19214,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(56));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_RNIIMEO9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(62),
cin => N_19213);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNILJA_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19212,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(55));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3_RNI067S8_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(63),
cin => N_19211);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIKIA_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19210,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(54));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3_RNIOAK3A_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(64),
cin => N_19209);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIJHA_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19208,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(53));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_RNICTUGA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(65),
cin => N_19207);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIIGA_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19206,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(52));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2_RNI92KV9_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(66),
cin => N_19205);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_RNIHFA_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19204,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(51));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1_RNIOH979_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1111000011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(67),
cin => N_19203);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD0_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19202,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.MIXOIN\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD0_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19201,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_U\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD0_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000010101010")
port map (
cout => N_19200,
dataa => VCC);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_REP1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_246_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(246),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(246));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_247_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100111101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(247),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(62),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(247));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_248_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100111101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(248),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(61),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(248));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_245_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(245),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(245),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_249_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(249),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(60),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(249),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\RETGRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_32_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => N_19149,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\RETGRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_SCTRL_NEW_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011000101")
port map (
combout => N_19148,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_A\(10));
\RETGRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_15_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => N_19147,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(49));
\RETGRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_15_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => N_19146,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_RNIBJRV_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_RNI9HRV_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPYBUS_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2_RETI\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_RNI7FRV_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_RNI5DRV_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(30));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_UN20_NOTSLRES: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES_RETI\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(31));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN13_NOTXZYFROMD_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1_RETI\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(49));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN13_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_RETI\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_RNIBNVV_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_RNIP3UV_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(49));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN13_NOTXZYFROMD_REP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2_RETI\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(49));
\GRLFPC20_R_FSR_CEXC_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1\(4),
dataa => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(4),
datab => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(4),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC20_R_FSR_CEXC_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1\(3),
dataa => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(3),
datab => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(3),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC20_R_FSR_CEXC_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1\(2),
dataa => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(2),
datab => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(2),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC20_R_FSR_CEXC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1\(1),
dataa => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(1),
datab => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(1),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC20_R_FSR_CEXC_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1\(0),
dataa => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(0),
datab => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(0),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(237),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(237),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(238),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(238),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(239),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(239),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(240),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(240),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(241),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(241),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(242),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(242),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(243),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(243),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(244),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(257),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(257),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(257),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(256),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(256),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(256),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(255),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(255),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(255),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(254),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(254),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(254),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(253),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(253),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(253),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(252),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(252),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(252),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(251),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(251),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(251),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(250),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(250),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(250),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\);
\GRLFPC20_R_I_RES_RNO_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.V.I.RES_1\(63),
dataa => \GRLFPC20.COMB.UN2_HOLDN\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT\,
datac => \GRLFPC20.COMB.V.I.RES_6_X\(63));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2S2_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_E\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN25_NOTXZYFROMD_RNIIJIB1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN15_NOTXZYFROMD_0_REP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN15_NOTXZYFROMD_0_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_XZBREGLOADEN_REP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_E\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN3_NOTXZYFROMD_RNIUMVM_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_WQSCTRL_RNILHL93_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN36_STKGEN_RNIJT6FH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010011111110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_S\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19_U\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN\);
\GRLFPC20_COMB_RS1_1_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.RS1_1_0_X\(3),
dataa => N_60,
datab => N_3,
datac => \GRLFPC20.R.A.RS1\(3));
\GRLFPC20_COMB_RS1_1_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.RS1_1_0_X\(4),
dataa => N_61,
datab => N_3,
datac => \GRLFPC20.R.A.RS1\(4));
\GRLFPC20_COMB_WRDATA_4_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(14),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(14),
datac => \GRLFPC20.R.I.RES\(43));
\GRLFPC20_COMB_WRDATA_4_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(46),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(46),
datac => \GRLFPC20.R.I.RES\(43));
\GRLFPC20_COMB_DBGDATA_4_0_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(10),
dataa => N_391,
datab => N_666,
datac => N_602);
\GRLFPC20_COMB_WRDATA_4_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(2),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(2),
datac => \GRLFPC20.R.I.RES\(31));
\GRLFPC20_COMB_WRDATA_4_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(11),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(11),
datac => \GRLFPC20.R.I.RES\(40));
\GRLFPC20_COMB_WRDATA_4_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(13),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(13),
datac => \GRLFPC20.R.I.RES\(42));
\GRLFPC20_COMB_WRDATA_4_X_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(17),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(17),
datac => \GRLFPC20.R.I.RES\(46));
\GRLFPC20_COMB_WRDATA_4_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(27),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(27),
datac => \GRLFPC20.R.I.RES\(56));
\GRLFPC20_COMB_WRDATA_4_X_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(29),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(29),
datac => \GRLFPC20.R.I.RES\(58));
\GRLFPC20_COMB_WRDATA_4_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(34),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(34),
datac => \GRLFPC20.R.I.RES\(31));
\GRLFPC20_COMB_WRDATA_4_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(43),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(43),
datac => \GRLFPC20.R.I.RES\(40));
\GRLFPC20_COMB_WRDATA_4_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(45),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(45),
datac => \GRLFPC20.R.I.RES\(42));
\GRLFPC20_COMB_WRDATA_4_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(49),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(49),
datac => \GRLFPC20.R.I.RES\(46));
\GRLFPC20_COMB_WRDATA_4_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(59),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(59),
datac => \GRLFPC20.R.I.RES\(56));
\GRLFPC20_COMB_WRDATA_4_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(61),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(61),
datac => \GRLFPC20.R.I.RES\(58));
\GRLFPC20_COMB_WRADDR_6_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.WRADDR_6_X\(3),
dataa => \GRLFPC20.WRADDR_1_SQMUXA\,
datab => N_347,
datac => \GRLFPC20.R.I.INST\(28));
\GRLFPC20_COMB_WRADDR_6_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.WRADDR_6_X\(4),
dataa => \GRLFPC20.WRADDR_1_SQMUXA\,
datab => N_348,
datac => \GRLFPC20.R.I.INST\(29));
\GRLFPC20_COMB_WRADDR_6_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.WRADDR_6_X\(1),
dataa => \GRLFPC20.WRADDR_1_SQMUXA\,
datab => N_345,
datac => \GRLFPC20.R.I.INST\(26));
\GRLFPC20_COMB_WRADDR_6_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.WRADDR_6_X\(2),
dataa => \GRLFPC20.WRADDR_1_SQMUXA\,
datab => N_346,
datac => \GRLFPC20.R.I.INST\(27));
\GRLFPC20_COMB_WRADDR_6_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.WRADDR_6_X\(0),
dataa => \GRLFPC20.WRADDR_1_SQMUXA\,
datab => N_344,
datac => \GRLFPC20.R.I.INST\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_102__G2_X\,
dataa => N_666,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_92__G2_X\,
dataa => N_676,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_COMB_DBGDATA_4_0_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(27),
dataa => N_391,
datab => N_683,
datac => N_619);
\GRLFPC20_COMB_WRDATA_4_X_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(21),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(21),
datac => \GRLFPC20.R.I.RES\(50));
\GRLFPC20_COMB_WRDATA_4_X_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(19),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(19),
datac => \GRLFPC20.R.I.RES\(48));
\GRLFPC20_COMB_WRDATA_4_X_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(18),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(18),
datac => \GRLFPC20.R.I.RES\(47));
\GRLFPC20_COMB_WRDATA_4_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(9),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(9),
datac => \GRLFPC20.R.I.RES\(38));
\GRLFPC20_COMB_WRDATA_4_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(38),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(38),
datac => \GRLFPC20.R.I.RES\(35));
\GRLFPC20_COMB_WRDATA_4_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(41),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(41),
datac => \GRLFPC20.R.I.RES\(38));
\GRLFPC20_COMB_WRDATA_4_X_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(12),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(12),
datac => \GRLFPC20.R.I.RES\(41));
\GRLFPC20_COMB_WRDATA_4_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(15),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(15),
datac => \GRLFPC20.R.I.RES\(44));
\GRLFPC20_COMB_WRDATA_4_X_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(20),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(20),
datac => \GRLFPC20.R.I.RES\(49));
\GRLFPC20_COMB_WRDATA_4_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(23),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(23),
datac => \GRLFPC20.R.I.RES\(52));
\GRLFPC20_COMB_WRDATA_4_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(44),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(44),
datac => \GRLFPC20.R.I.RES\(41));
\GRLFPC20_COMB_WRDATA_4_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(47),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(47),
datac => \GRLFPC20.R.I.RES\(44));
\GRLFPC20_COMB_WRDATA_4_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(52),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(52),
datac => \GRLFPC20.R.I.RES\(49));
\GRLFPC20_COMB_WRDATA_4_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(55),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(55),
datac => \GRLFPC20.R.I.RES\(52));
\GRLFPC20_FPI_OP1_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(44),
dataa => N_668,
datab => N_604,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(47),
dataa => N_671,
datab => N_607,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_DBGDATA_4_0_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(7),
dataa => N_391,
datab => N_663,
datac => N_599);
\GRLFPC20_COMB_DBGDATA_4_0_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(15),
dataa => N_391,
datab => N_671,
datac => N_607);
\GRLFPC20_COMB_V_FSR_FCC_1_1_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC_1_1_X\(0),
dataa => N_366,
datab => CPO_CCZ(0),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_COMB_V_FSR_FCC_1_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC_1_1_X\(1),
dataa => N_367,
datab => CPO_CCZ(1),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_105__G2_X\,
dataa => N_663,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_103__G2_X\,
dataa => N_665,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_100__G2_X\,
dataa => N_668,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_97__G2_X\,
dataa => N_671,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_COMB_DBGDATA_4_0_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(9),
dataa => N_391,
datab => N_665,
datac => N_601);
\GRLFPC20_COMB_WRDATA_4_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(50),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(50),
datac => \GRLFPC20.R.I.RES\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_99__G2_X\,
dataa => N_669,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_COMB_DBGDATA_4_0_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(13),
dataa => N_391,
datab => N_669,
datac => N_605);
GRLFPC20_COMB_FPDECODE_FPOP2_0_O2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC20.COMB.FPDECODE.FPOP2_0_O2_X\,
dataa => N_67,
datab => N_65);
GRLFPC20_COMB_FPDECODE_FPOP8_I_O3_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC20.COMB.FPDECODE.FPOP8_I_O3_X\,
dataa => N_74,
datab => N_73);
GRLFPC20_RS2_0_SQMUXA_RNI7CQD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.COMB.RS1_1_SN_M2_X\,
dataa => N_3,
datab => \GRLFPC20.RS2_0_SQMUXA\);
GRLFPC20_COMB_V_A_RF1REN_1_0_650_A2_3_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.COMB.V.A.RF1REN_1_0_650_A2_3_X\,
dataa => N_73,
datab => N_74);
\GRLFPC20_COMB_WRDATA_4_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(8),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(8),
datac => \GRLFPC20.R.I.RES\(37));
\GRLFPC20_COMB_WRDATA_4_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(40),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(40),
datac => \GRLFPC20.R.I.RES\(37));
\GRLFPC20_COMB_DBGDATA_4_0_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(23),
dataa => N_391,
datab => N_679,
datac => N_615);
\GRLFPC20_COMB_DBGDATA_4_0_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(25),
dataa => N_391,
datab => N_681,
datac => N_617);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_89__G2_X\,
dataa => N_679,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
GRLFPC20_COMB_UN3_HOLDN_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.COMB.UN3_HOLDN_X\,
dataa => N_146,
datab => N_147);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_84__G2_X\,
dataa => N_684,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_87__G2_X\,
dataa => N_681,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_FPI_OP1_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(60),
dataa => N_684,
datab => N_620,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
GRLFPC20_COMB_V_E_STDATA2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA2_X\,
dataa => N_145,
datab => N_144);
GRLFPC20_COMB_RSDECODE_RS1V_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.COMB.RSDECODE.RS1V_X\,
dataa => N_76,
datab => N_75);
GRLFPC20_R_MK_HOLDN1_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC20.R.MK.HOLDN1_0_0_G0_X\,
dataa => N_1,
datab => \GRLFPC20.R.MK.RST2\);
\GRLFPC20_FPI_OP1_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(63),
dataa => N_687,
datab => N_623,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP2_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(63),
dataa => N_719,
datab => N_655,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_COMB_WRDATA_4_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(7),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(7),
datac => \GRLFPC20.R.I.RES\(36));
\GRLFPC20_COMB_WRDATA_4_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(10),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(10),
datac => \GRLFPC20.R.I.RES\(39));
\GRLFPC20_COMB_WRDATA_4_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(24),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(24),
datac => \GRLFPC20.R.I.RES\(53));
\GRLFPC20_COMB_WRDATA_4_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(31),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(31),
datac => \GRLFPC20.R.I.RES\(63));
\GRLFPC20_COMB_WRDATA_4_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(36),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(36),
datac => \GRLFPC20.R.I.RES\(33));
\GRLFPC20_COMB_WRDATA_4_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(39),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(39),
datac => \GRLFPC20.R.I.RES\(36));
\GRLFPC20_COMB_WRDATA_4_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(42),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(42),
datac => \GRLFPC20.R.I.RES\(39));
\GRLFPC20_COMB_WRDATA_4_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(56),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(56),
datac => \GRLFPC20.R.I.RES\(53));
\GRLFPC20_FPI_OP1_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(38),
dataa => N_662,
datab => N_598,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_DBGDATA_4_0_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(6),
dataa => N_391,
datab => N_662,
datac => N_598);
\GRLFPC20_COMB_DBGDATA_4_0_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(24),
dataa => N_391,
datab => N_680,
datac => N_616);
\GRLFPC20_WRDATA_0_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(63),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_387,
datac => \GRLFPC20.R.I.RES\(63));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_85__G2_X\,
dataa => N_683,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_COMB_WRDATA_4_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(62),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(62),
datac => \GRLFPC20.R.I.RES\(59));
\GRLFPC20_COMB_WRDATA_4_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(33),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(33),
datac => \GRLFPC20.R.I.RES\(30));
\GRLFPC20_COMB_WRDATA_4_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(30),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(30),
datac => \GRLFPC20.R.I.RES\(59));
\GRLFPC20_COMB_WRDATA_4_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(60),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(60),
datac => \GRLFPC20.R.I.RES\(57));
\GRLFPC20_COMB_WRDATA_4_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(53),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(53),
datac => \GRLFPC20.R.I.RES\(50));
\GRLFPC20_COMB_WRDATA_4_X_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(28),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(28),
datac => \GRLFPC20.R.I.RES\(57));
\GRLFPC20_COMB_WRDATA_4_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(22),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(22),
datac => \GRLFPC20.R.I.RES\(51));
\GRLFPC20_COMB_WRDATA_4_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(51),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(51),
datac => \GRLFPC20.R.I.RES\(48));
\GRLFPC20_COMB_WRDATA_4_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(54),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(54),
datac => \GRLFPC20.R.I.RES\(51));
\GRLFPC20_FPI_OP1_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(51),
dataa => N_675,
datab => N_611,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(54),
dataa => N_678,
datab => N_614,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(57),
dataa => N_681,
datab => N_617,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_DBGDATA_4_0_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(22),
dataa => N_391,
datab => N_678,
datac => N_614);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_90__G2_X\,
dataa => N_678,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_FPI_OP1_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(59),
dataa => N_683,
datab => N_619,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(62),
dataa => N_686,
datab => N_622,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_DBGDATA_4_0_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(30),
dataa => N_391,
datab => N_686,
datac => N_622);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_108__G2_X\,
dataa => N_660,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
GRLFPC20_COMB_RDD_1_M10_2_0_A2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.COMB.RDD_1.M10_2_0_A2_X\,
dataa => N_63,
datab => N_62);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_MAPMULXFF_UN4_UNIMPMAP_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_1_X\,
dataa => N_52,
datab => N_55);
\GRLFPC20_COMB_WRDATA_4_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(0),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(0),
datac => \GRLFPC20.R.I.RES\(29));
\GRLFPC20_COMB_WRDATA_4_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(1),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(1),
datac => \GRLFPC20.R.I.RES\(30));
\GRLFPC20_COMB_WRDATA_4_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(5),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(5),
datac => \GRLFPC20.R.I.RES\(34));
\GRLFPC20_COMB_DBGDATA_4_0_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(5),
dataa => N_391,
datab => N_661,
datac => N_597);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_107__G2_X\,
dataa => N_661,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
GRLFPC20_RS1D_CNST_0_A2_2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.RS1D_CNST_0_A2_2_X\,
dataa => N_67,
datab => N_64);
\GRLFPC20_COMB_RS1_1_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.RS1_1_0_X\(2),
dataa => N_59,
datab => N_3,
datac => \GRLFPC20.R.A.RS1\(2));
\GRLFPC20_COMB_RS1_1_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.RS1_1_0_X\(0),
dataa => N_57,
datab => N_3,
datac => \GRLFPC20.R.A.RS1\(0));
\GRLFPC20_FPI_OP1_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(45),
dataa => N_669,
datab => N_605,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_DBGDATA_4_0_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(16),
dataa => N_391,
datab => N_672,
datac => N_608);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_96__G2_X\,
dataa => N_672,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_COMB_DBGDATA_4_0_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(31),
dataa => N_391,
datab => N_687,
datac => N_623);
\GRLFPC20_R_FSR_TEM_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.TEM_1_0_4__G3_X\,
dataa => N_383,
datab => \GRLFPC20.R.FSR.TEM\(4),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_R_FSR_TEM_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.TEM_1_0_3__G3_X\,
dataa => N_382,
datab => \GRLFPC20.R.FSR.TEM\(3),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_R_FSR_TEM_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.TEM_1_0_2__G3_X\,
dataa => N_381,
datab => \GRLFPC20.R.FSR.TEM\(2),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_R_FSR_TEM_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.TEM_1_0_1__G3_X\,
dataa => N_380,
datab => \GRLFPC20.R.FSR.TEM\(1),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_R_FSR_TEM_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.TEM_1_0_0__G3_X\,
dataa => N_379,
datab => \GRLFPC20.R.FSR.TEM\(0),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_R_FSR_RD_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.RD_0_0_1__G3_X\,
dataa => N_387,
datab => \GRLFPC20.R.FSR.RD\(1),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_R_FSR_RD_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.RD_0_0_0__G3_X\,
dataa => N_386,
datab => \GRLFPC20.R.FSR.RD\(0),
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
GRLFPC20_R_FSR_NONSTD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.R.FSR.NONSTD_0_0_G3_X\,
dataa => N_378,
datab => \GRLFPC20.R.FSR.NONSTD\,
datac => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_86__G2_X\,
dataa => N_682,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_88__G2_X\,
dataa => N_680,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_91__G2_X\,
dataa => N_677,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_93__G2_X\,
dataa => N_675,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_94__G2_X\,
dataa => N_674,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_95__G2_X\,
dataa => N_673,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_98__G2_X\,
dataa => N_670,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_101__G2_X\,
dataa => N_667,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_104__G2_X\,
dataa => N_664,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_106__G2_X\,
dataa => N_662,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_109__G2_X\,
dataa => N_659,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_110__G2_X\,
dataa => N_658,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_111__G2_X\,
dataa => N_657,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_112__G2_X\,
dataa => N_656,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11));
\GRLFPC20_FPI_OP2_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(32),
dataa => N_688,
datab => N_624,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(33),
dataa => N_689,
datab => N_625,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(34),
dataa => N_690,
datab => N_626,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(35),
dataa => N_691,
datab => N_627,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(36),
dataa => N_692,
datab => N_628,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(37),
dataa => N_693,
datab => N_629,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(38),
dataa => N_694,
datab => N_630,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(39),
dataa => N_695,
datab => N_631,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(40),
dataa => N_696,
datab => N_632,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(41),
dataa => N_697,
datab => N_633,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(42),
dataa => N_698,
datab => N_634,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(43),
dataa => N_699,
datab => N_635,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(44),
dataa => N_700,
datab => N_636,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(45),
dataa => N_701,
datab => N_637,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(46),
dataa => N_702,
datab => N_638,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(47),
dataa => N_703,
datab => N_639,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(48),
dataa => N_704,
datab => N_640,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(49),
dataa => N_705,
datab => N_641,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(50),
dataa => N_706,
datab => N_642,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(51),
dataa => N_707,
datab => N_643,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(52),
dataa => N_708,
datab => N_644,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(53),
dataa => N_709,
datab => N_645,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(54),
dataa => N_710,
datab => N_646,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(55),
dataa => N_711,
datab => N_647,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(56),
dataa => N_712,
datab => N_648,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(57),
dataa => N_713,
datab => N_649,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(58),
dataa => N_714,
datab => N_650,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(59),
dataa => N_715,
datab => N_651,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(60),
dataa => N_716,
datab => N_652,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(61),
dataa => N_717,
datab => N_653,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP2_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP2_X\(62),
dataa => N_718,
datab => N_654,
datac => \GRLFPC20.COMB.UN1_FPCI_4\);
\GRLFPC20_FPI_OP1_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(35),
dataa => N_659,
datab => N_595,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(41),
dataa => N_665,
datab => N_601,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_DBGDATA_4_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(3),
dataa => N_391,
datab => N_659,
datac => N_595);
\GRLFPC20_COMB_WRDATA_4_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(58),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(58),
datac => \GRLFPC20.R.I.RES\(55));
\GRLFPC20_COMB_WRDATA_4_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(26),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(26),
datac => \GRLFPC20.R.I.RES\(55));
\GRLFPC20_COMB_V_FSR_CEXC_1_1_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(4),
dataa => N_360,
datab => \GRLFPC20.R.FSR.CEXC\(4),
datac => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC20_COMB_V_FSR_CEXC_1_1_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(3),
dataa => N_359,
datab => \GRLFPC20.R.FSR.CEXC\(3),
datac => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC20_COMB_V_FSR_CEXC_1_1_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(2),
dataa => N_358,
datab => \GRLFPC20.R.FSR.CEXC\(2),
datac => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC20_COMB_V_FSR_CEXC_1_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(1),
dataa => N_357,
datab => \GRLFPC20.R.FSR.CEXC\(1),
datac => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC20_COMB_V_FSR_CEXC_1_1_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_1_X\(0),
dataa => N_356,
datab => \GRLFPC20.R.FSR.CEXC\(0),
datac => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC20_COMB_DBGDATA_4_0_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(26),
dataa => N_391,
datab => N_682,
datac => N_618);
\GRLFPC20_COMB_DBGDATA_4_0_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(14),
dataa => N_391,
datab => N_670,
datac => N_606);
\GRLFPC20_COMB_DBGDATA_4_0_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(11),
dataa => N_391,
datab => N_667,
datac => N_603);
\GRLFPC20_COMB_DBGDATA_4_0_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(8),
dataa => N_391,
datab => N_664,
datac => N_600);
\GRLFPC20_COMB_DBGDATA_4_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(4),
dataa => N_391,
datab => N_660,
datac => N_596);
\GRLFPC20_COMB_DBGDATA_4_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(2),
dataa => N_391,
datab => N_658,
datac => N_594);
\GRLFPC20_COMB_DBGDATA_4_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(1),
dataa => N_391,
datab => N_657,
datac => N_593);
\GRLFPC20_COMB_DBGDATA_4_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.DBGDATA_4_0_X\(0),
dataa => N_391,
datab => N_656,
datac => N_592);
\GRLFPC20_FPI_OP1_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(58),
dataa => N_682,
datab => N_618,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(56),
dataa => N_680,
datab => N_616,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(55),
dataa => N_679,
datab => N_615,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(53),
dataa => N_677,
datab => N_613,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(52),
dataa => N_676,
datab => N_612,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(50),
dataa => N_674,
datab => N_610,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(49),
dataa => N_673,
datab => N_609,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(48),
dataa => N_672,
datab => N_608,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(46),
dataa => N_670,
datab => N_606,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(43),
dataa => N_667,
datab => N_603,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(42),
dataa => N_666,
datab => N_602,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(40),
dataa => N_664,
datab => N_600,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(39),
dataa => N_663,
datab => N_599,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(37),
dataa => N_661,
datab => N_597,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(36),
dataa => N_660,
datab => N_596,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(34),
dataa => N_658,
datab => N_594,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(33),
dataa => N_657,
datab => N_593,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_FPI_OP1_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(32),
dataa => N_656,
datab => N_592,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_WRDATA_4_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(57),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(57),
datac => \GRLFPC20.R.I.RES\(54));
\GRLFPC20_COMB_WRDATA_4_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(37),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(37),
datac => \GRLFPC20.R.I.RES\(34));
\GRLFPC20_COMB_WRDATA_4_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(32),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(32),
datac => \GRLFPC20.R.I.RES\(29));
\GRLFPC20_COMB_WRDATA_4_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(25),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(25),
datac => \GRLFPC20.R.I.RES\(54));
\GRLFPC20_COMB_WRDATA_4_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(4),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(4),
datac => \GRLFPC20.R.I.RES\(33));
\GRLFPC20_FPI_OP1_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.FPI.OP1_X\(61),
dataa => N_685,
datab => N_621,
datac => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_COMB_WRDATA_4_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(48),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(48),
datac => \GRLFPC20.R.I.RES\(45));
\GRLFPC20_COMB_WRDATA_4_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(35),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(35),
datac => \GRLFPC20.R.I.RES\(32));
\GRLFPC20_COMB_WRDATA_4_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(16),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(16),
datac => \GRLFPC20.R.I.RES\(45));
\GRLFPC20_COMB_WRDATA_4_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(6),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(6),
datac => \GRLFPC20.R.I.RES\(35));
\GRLFPC20_COMB_WRDATA_4_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.WRDATA_4_X\(3),
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.R.I.RES\(3),
datac => \GRLFPC20.R.I.RES\(32));
\GRLFPC20_COMB_RS1_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.RS1_1_0_X\(1),
dataa => N_58,
datab => N_3,
datac => \GRLFPC20.R.A.RS1\(1));
GRLFPC20_COMB_FPDECODE_RDD5_3_0_A2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.COMB.FPDECODE.RDD5_3_0_A2_X\,
dataa => N_53,
datab => N_52);
GRLFPC20_R_I_V_RNIKG6C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_0_X\,
dataa => N_1,
datab => \GRLFPC20.R.I.V\);
GRLFPC20_COMB_LOCK_1_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.COMB.LOCK_1_1_X\,
dataa => N_78,
datab => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\);
GRLFPC20_RS1D_CNST_0_A2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.RS1D_CNST_0_A2_1_X\,
dataa => N_65,
datab => N_74);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_0__G0_0_A3_0_X\,
dataa => N_55,
datab => N_51);
GRLFPC20_COMB_UN1_FPCI_4_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.COMB.UN1_FPCI_0_1_X\,
dataa => N_145,
datab => \GRLFPC20.R.A.ST\);
GRLFPC20_WREN1_0_SQMUXA_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.WREN1_0_SQMUXA_1_X\,
dataa => N_339,
datab => \GRLFPC20.R.X.AFSR\,
datac => \GRLFPC20.R.X.LD\);
\GRLFPC20_COMB_DBGDATA_4_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(10),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(10),
datac => CPO_CCZ(0));
\GRLFPC20_WRDATA_0_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(14),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_370,
datac => \GRLFPC20.COMB.WRDATA_4_X\(14));
\GRLFPC20_WRDATA_0_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(46),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_370,
datac => \GRLFPC20.COMB.WRDATA_4_X\(46));
\GRLFPC20_WRDATA_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(2),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_358,
datac => \GRLFPC20.COMB.WRDATA_4_X\(2));
\GRLFPC20_WRDATA_0_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(11),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_367,
datac => \GRLFPC20.COMB.WRDATA_4_X\(11));
\GRLFPC20_WRDATA_0_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(13),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_369,
datac => \GRLFPC20.COMB.WRDATA_4_X\(13));
\GRLFPC20_WRDATA_0_X_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(17),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_373,
datac => \GRLFPC20.COMB.WRDATA_4_X\(17));
\GRLFPC20_WRDATA_0_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(27),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_383,
datac => \GRLFPC20.COMB.WRDATA_4_X\(27));
\GRLFPC20_WRDATA_0_X_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(29),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_385,
datac => \GRLFPC20.COMB.WRDATA_4_X\(29));
\GRLFPC20_WRDATA_0_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(34),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_358,
datac => \GRLFPC20.COMB.WRDATA_4_X\(34));
\GRLFPC20_WRDATA_0_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(43),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_367,
datac => \GRLFPC20.COMB.WRDATA_4_X\(43));
\GRLFPC20_WRDATA_0_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(45),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_369,
datac => \GRLFPC20.COMB.WRDATA_4_X\(45));
\GRLFPC20_WRDATA_0_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(49),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_373,
datac => \GRLFPC20.COMB.WRDATA_4_X\(49));
\GRLFPC20_WRDATA_0_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(59),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_383,
datac => \GRLFPC20.COMB.WRDATA_4_X\(59));
\GRLFPC20_WRDATA_0_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(61),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_385,
datac => \GRLFPC20.COMB.WRDATA_4_X\(61));
\GRLFPC20_COMB_DBGDATA_4_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(27),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(27),
datac => \GRLFPC20.R.FSR.TEM\(4));
\GRLFPC20_WRDATA_0_X_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(21),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_377,
datac => \GRLFPC20.COMB.WRDATA_4_X\(21));
\GRLFPC20_WRDATA_0_X_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(19),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_375,
datac => \GRLFPC20.COMB.WRDATA_4_X\(19));
\GRLFPC20_WRDATA_0_X_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(18),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_374,
datac => \GRLFPC20.COMB.WRDATA_4_X\(18));
\GRLFPC20_WRDATA_0_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(9),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_365,
datac => \GRLFPC20.COMB.WRDATA_4_X\(9));
\GRLFPC20_WRDATA_0_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(38),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_362,
datac => \GRLFPC20.COMB.WRDATA_4_X\(38));
\GRLFPC20_WRDATA_0_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(41),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_365,
datac => \GRLFPC20.COMB.WRDATA_4_X\(41));
\GRLFPC20_COMB_DBGDATA_4_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(7),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(7),
datac => \GRLFPC20.R.FSR.AEXC\(2));
\GRLFPC20_COMB_DBGDATA_4_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(15),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(15),
datac => \GRLFPC20.R.FSR.FTT\(1));
\GRLFPC20_WRDATA_0_X_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(12),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_368,
datac => \GRLFPC20.COMB.WRDATA_4_X\(12));
\GRLFPC20_WRDATA_0_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(15),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_371,
datac => \GRLFPC20.COMB.WRDATA_4_X\(15));
\GRLFPC20_WRDATA_0_X_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(20),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_376,
datac => \GRLFPC20.COMB.WRDATA_4_X\(20));
\GRLFPC20_WRDATA_0_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(23),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_379,
datac => \GRLFPC20.COMB.WRDATA_4_X\(23));
\GRLFPC20_WRDATA_0_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(44),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_368,
datac => \GRLFPC20.COMB.WRDATA_4_X\(44));
\GRLFPC20_WRDATA_0_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(47),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_371,
datac => \GRLFPC20.COMB.WRDATA_4_X\(47));
\GRLFPC20_WRDATA_0_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(52),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_376,
datac => \GRLFPC20.COMB.WRDATA_4_X\(52));
\GRLFPC20_WRDATA_0_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(55),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_379,
datac => \GRLFPC20.COMB.WRDATA_4_X\(55));
\GRLFPC20_COMB_DBGDATA_4_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(9),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(9),
datac => \GRLFPC20.R.FSR.AEXC\(4));
\GRLFPC20_WRDATA_0_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(50),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_374,
datac => \GRLFPC20.COMB.WRDATA_4_X\(50));
GRLFPC20_WRADDR_0_SQMUXA_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.WRADDR_0_SQMUXA_X\,
dataa => N_390,
datab => N_389,
datac => N_388);
\GRLFPC20_COMB_DBGDATA_4_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(23),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(23),
datac => \GRLFPC20.R.FSR.TEM\(0));
\GRLFPC20_COMB_DBGDATA_4_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(25),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(25),
datac => \GRLFPC20.R.FSR.TEM\(2));
\GRLFPC20_WRDATA_0_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(8),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_364,
datac => \GRLFPC20.COMB.WRDATA_4_X\(8));
\GRLFPC20_WRDATA_0_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(40),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_364,
datac => \GRLFPC20.COMB.WRDATA_4_X\(40));
GRLFPC20_R_E_AFQ_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.E.AFQ_0_0_G1_X\,
dataa => N_147,
datab => N_146,
datac => \GRLFPC20.R.A.AFQ\);
GRLFPC20_R_E_AFSR_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.E.AFSR_0_0_G1_X\,
dataa => N_147,
datab => N_146,
datac => \GRLFPC20.R.A.AFSR\);
GRLFPC20_R_E_FPOP_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.E.FPOP_0_0_G1_X\,
dataa => N_147,
datab => N_146,
datac => \GRLFPC20.R.A.FPOP\);
GRLFPC20_R_E_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.E.LD_0_0_G1_X\,
dataa => N_147,
datab => N_146,
datac => \GRLFPC20.R.A.LD\);
GRLFPC20_ANNULFPU_0_SQMUXA_2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000011100000")
port map (
combout => \GRLFPC20.ANNULFPU_0_SQMUXA_2_X\,
dataa => N_147,
datab => N_146,
datac => \GRLFPC20.R.A.FPOP\);
\GRLFPC20_COMB_V_E_STDATA_1_0_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(27),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(27),
datac => \GRLFPC20.R.I.INST\(27));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(26),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(26),
datac => \GRLFPC20.R.I.INST\(26));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(25),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(25),
datac => \GRLFPC20.R.I.INST\(25));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(31),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(31),
datac => \GRLFPC20.R.I.INST\(31));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(30),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(30),
datac => \GRLFPC20.R.I.INST\(30));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(24),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(24),
datac => \GRLFPC20.R.I.INST\(24));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(23),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(23),
datac => \GRLFPC20.R.I.INST\(23));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(22),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(22),
datac => \GRLFPC20.R.I.INST\(22));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(16),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(16),
datac => \GRLFPC20.R.I.INST\(16));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(15),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(15),
datac => \GRLFPC20.R.I.INST\(15));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(14),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(14),
datac => \GRLFPC20.R.I.INST\(14));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(13),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(13),
datac => \GRLFPC20.R.I.INST\(13));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(11),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(11),
datac => \GRLFPC20.R.I.INST\(11));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(10),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(10),
datac => \GRLFPC20.R.I.INST\(10));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(9),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(9),
datac => \GRLFPC20.R.I.INST\(9));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(8),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(8),
datac => \GRLFPC20.R.I.INST\(8));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(7),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(7),
datac => \GRLFPC20.R.I.INST\(7));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(6),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(6),
datac => \GRLFPC20.R.I.INST\(6));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(5),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(5),
datac => \GRLFPC20.R.I.INST\(5));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(4),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(4),
datac => \GRLFPC20.R.I.INST\(4));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(3),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(3),
datac => \GRLFPC20.R.I.INST\(3));
\GRLFPC20_COMB_V_E_STDATA_1_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(2),
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(2),
datac => \GRLFPC20.R.I.INST\(2));
\GRLFPC20_R_E_STDATA_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000011010000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_0__G3_X\,
dataa => N_144,
datab => N_145,
datac => \GRLFPC20.R.I.INST\(0));
\GRLFPC20_R_E_STDATA_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000011010000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_1__G3_X\,
dataa => N_144,
datab => N_145,
datac => \GRLFPC20.R.I.INST\(1));
\GRLFPC20_R_E_STDATA_RNO_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_12__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(12),
datac => \GRLFPC20.R.I.INST\(12));
\GRLFPC20_R_E_STDATA_RNO_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_17__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(17),
datac => \GRLFPC20.R.I.INST\(17));
\GRLFPC20_R_E_STDATA_RNO_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_18__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(18),
datac => \GRLFPC20.R.I.INST\(18));
\GRLFPC20_R_E_STDATA_RNO_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_19__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(19),
datac => \GRLFPC20.R.I.INST\(19));
\GRLFPC20_R_E_STDATA_RNO_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_20__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(20),
datac => \GRLFPC20.R.I.INST\(20));
\GRLFPC20_R_E_STDATA_RNO_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_21__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(21),
datac => \GRLFPC20.R.I.INST\(21));
\GRLFPC20_R_E_STDATA_RNO_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_28__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(28),
datac => \GRLFPC20.R.I.INST\(28));
\GRLFPC20_R_E_STDATA_RNO_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_29__G3_X\,
dataa => \GRLFPC20.COMB.V.E.STDATA2_X\,
datab => \GRLFPC20.R.I.PC\(29),
datac => \GRLFPC20.R.I.INST\(29));
GRLFPC20_R_M_AFQ_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.M.AFQ_0_0_G1_X\,
dataa => N_216,
datab => N_215,
datac => \GRLFPC20.R.E.AFQ\);
GRLFPC20_R_M_AFSR_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.M.AFSR_0_0_G1_X\,
dataa => N_216,
datab => N_215,
datac => \GRLFPC20.R.E.AFSR\);
GRLFPC20_R_M_FPOP_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.M.FPOP_0_0_G1_X\,
dataa => N_216,
datab => N_215,
datac => \GRLFPC20.R.E.FPOP\);
GRLFPC20_R_M_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.M.LD_0_0_G1_X\,
dataa => N_216,
datab => N_215,
datac => \GRLFPC20.R.E.LD\);
GRLFPC20_R_X_AFQ_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.X.AFQ_0_0_G1_X\,
dataa => N_285,
datab => N_284,
datac => \GRLFPC20.R.M.AFQ\);
GRLFPC20_R_X_AFSR_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.X.AFSR_0_0_G1_X\,
dataa => N_285,
datab => N_284,
datac => \GRLFPC20.R.M.AFSR\);
GRLFPC20_R_X_FPOP_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.X.FPOP_0_0_G1_X\,
dataa => N_285,
datab => N_284,
datac => \GRLFPC20.R.M.FPOP\);
GRLFPC20_R_X_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.R.X.LD_0_0_G1_X\,
dataa => N_285,
datab => N_284,
datac => \GRLFPC20.R.M.LD\);
GRLFPC20_ANNULFPU_0_SQMUXA_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000011100000")
port map (
combout => \GRLFPC20.ANNULFPU_0_SQMUXA_1_X\,
dataa => N_216,
datab => N_215,
datac => \GRLFPC20.R.E.FPOP\);
GRLFPC20_ANNULFPU_0_SQMUXA_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000011100000")
port map (
combout => \GRLFPC20.ANNULFPU_0_SQMUXA_X\,
dataa => N_285,
datab => N_284,
datac => \GRLFPC20.R.M.FPOP\);
\GRLFPC20_COMB_DBGDATA_4_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(6),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(6),
datac => \GRLFPC20.R.FSR.AEXC\(1));
\GRLFPC20_COMB_DBGDATA_4_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(24),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(24),
datac => \GRLFPC20.R.FSR.TEM\(1));
\GRLFPC20_WRDATA_0_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(7),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_363,
datac => \GRLFPC20.COMB.WRDATA_4_X\(7));
\GRLFPC20_WRDATA_0_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(10),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_366,
datac => \GRLFPC20.COMB.WRDATA_4_X\(10));
\GRLFPC20_WRDATA_0_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(24),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_380,
datac => \GRLFPC20.COMB.WRDATA_4_X\(24));
\GRLFPC20_WRDATA_0_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(31),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_387,
datac => \GRLFPC20.COMB.WRDATA_4_X\(31));
\GRLFPC20_WRDATA_0_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(36),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_360,
datac => \GRLFPC20.COMB.WRDATA_4_X\(36));
\GRLFPC20_WRDATA_0_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(39),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_363,
datac => \GRLFPC20.COMB.WRDATA_4_X\(39));
\GRLFPC20_WRDATA_0_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(42),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_366,
datac => \GRLFPC20.COMB.WRDATA_4_X\(42));
\GRLFPC20_WRDATA_0_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(56),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_380,
datac => \GRLFPC20.COMB.WRDATA_4_X\(56));
\GRLFPC20_WRDATA_0_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(62),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_386,
datac => \GRLFPC20.COMB.WRDATA_4_X\(62));
\GRLFPC20_WRDATA_0_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(33),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_357,
datac => \GRLFPC20.COMB.WRDATA_4_X\(33));
\GRLFPC20_WRDATA_0_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(30),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_386,
datac => \GRLFPC20.COMB.WRDATA_4_X\(30));
\GRLFPC20_WRDATA_0_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(60),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_384,
datac => \GRLFPC20.COMB.WRDATA_4_X\(60));
\GRLFPC20_WRDATA_0_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(53),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_377,
datac => \GRLFPC20.COMB.WRDATA_4_X\(53));
\GRLFPC20_WRDATA_0_X_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(28),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_384,
datac => \GRLFPC20.COMB.WRDATA_4_X\(28));
\GRLFPC20_WRDATA_0_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(22),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_378,
datac => \GRLFPC20.COMB.WRDATA_4_X\(22));
\GRLFPC20_COMB_DBGDATA_4_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(22),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(22),
datac => \GRLFPC20.R.FSR.NONSTD\);
\GRLFPC20_WRDATA_0_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(51),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_375,
datac => \GRLFPC20.COMB.WRDATA_4_X\(51));
\GRLFPC20_WRDATA_0_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(54),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_378,
datac => \GRLFPC20.COMB.WRDATA_4_X\(54));
\GRLFPC20_COMB_DBGDATA_4_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(30),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(30),
datac => \GRLFPC20.R.FSR.RD\(0));
\GRLFPC20_COMB_DBGDATA_4_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(5),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(5),
datac => \GRLFPC20.R.FSR.AEXC\(0));
\GRLFPC20_WRDATA_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(0),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_356,
datac => \GRLFPC20.COMB.WRDATA_4_X\(0));
\GRLFPC20_WRDATA_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(1),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_357,
datac => \GRLFPC20.COMB.WRDATA_4_X\(1));
\GRLFPC20_WRDATA_0_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(5),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_361,
datac => \GRLFPC20.COMB.WRDATA_4_X\(5));
GRLFPC20_COMB_FPDECODE_RDD4_0_A2_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.RDD4_0_A2_0_X\,
dataa => N_51,
datab => N_50,
datac => N_53);
\GRLFPC20_COMB_DBGDATA_4_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(16),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(16),
datac => \GRLFPC20.R.FSR.FTT\(2));
\GRLFPC20_COMB_DBGDATA_4_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(31),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(31),
datac => \GRLFPC20.R.FSR.RD\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1_X\(23),
dataa => N_719,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP2_X\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1_X\(25),
dataa => N_717,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP2_X\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1_X\(24),
dataa => N_718,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP2_X\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_X_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_X\(81),
dataa => N_687,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP1_X\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_X_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_X\(83),
dataa => N_685,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP1_X\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_X_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_X\(82),
dataa => N_686,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP1_X\(33));
\GRLFPC20_WRDATA_0_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(58),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_382,
datac => \GRLFPC20.COMB.WRDATA_4_X\(58));
\GRLFPC20_WRDATA_0_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(26),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_382,
datac => \GRLFPC20.COMB.WRDATA_4_X\(26));
\GRLFPC20_COMB_DBGDATA_4_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(3),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(3),
datac => \GRLFPC20.R.FSR.CEXC\(3));
\GRLFPC20_WRDATA_0_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(57),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_381,
datac => \GRLFPC20.COMB.WRDATA_4_X\(57));
\GRLFPC20_WRDATA_0_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(37),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_361,
datac => \GRLFPC20.COMB.WRDATA_4_X\(37));
\GRLFPC20_WRDATA_0_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(32),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_356,
datac => \GRLFPC20.COMB.WRDATA_4_X\(32));
\GRLFPC20_WRDATA_0_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(25),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_381,
datac => \GRLFPC20.COMB.WRDATA_4_X\(25));
\GRLFPC20_WRDATA_0_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(4),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_360,
datac => \GRLFPC20.COMB.WRDATA_4_X\(4));
\GRLFPC20_COMB_DBGDATA_4_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(26),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(26),
datac => \GRLFPC20.R.FSR.TEM\(3));
\GRLFPC20_COMB_DBGDATA_4_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(14),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(14),
datac => \GRLFPC20.R.FSR.FTT\(0));
\GRLFPC20_COMB_DBGDATA_4_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(11),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(11),
datac => CPO_CCZ(1));
\GRLFPC20_COMB_DBGDATA_4_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(8),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(8),
datac => \GRLFPC20.R.FSR.AEXC\(3));
\GRLFPC20_COMB_DBGDATA_4_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(4),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(4),
datac => \GRLFPC20.R.FSR.CEXC\(4));
\GRLFPC20_COMB_DBGDATA_4_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(2),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(2),
datac => \GRLFPC20.R.FSR.CEXC\(2));
\GRLFPC20_COMB_DBGDATA_4_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(1),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(1),
datac => \GRLFPC20.R.FSR.CEXC\(1));
\GRLFPC20_COMB_DBGDATA_4_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => CPO_DBG_DATAZ(0),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(0),
datac => \GRLFPC20.R.FSR.CEXC\(0));
\GRLFPC20_WRDATA_0_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(48),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_372,
datac => \GRLFPC20.COMB.WRDATA_4_X\(48));
\GRLFPC20_WRDATA_0_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(35),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_359,
datac => \GRLFPC20.COMB.WRDATA_4_X\(35));
\GRLFPC20_WRDATA_0_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(16),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_372,
datac => \GRLFPC20.COMB.WRDATA_4_X\(16));
\GRLFPC20_WRDATA_0_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(6),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_362,
datac => \GRLFPC20.COMB.WRDATA_4_X\(6));
\GRLFPC20_WRDATA_0_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.WRDATA_0_X\(3),
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => N_359,
datac => \GRLFPC20.COMB.WRDATA_4_X\(3));
GRLFPC20_COMB_FPDECODE_RDD4_0_A2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.COMB.FPDECODE.RDD4_0_A2_X\,
dataa => N_49,
datab => N_48,
datac => N_54);
GRLFPC20_COMB_RSDECODE_UN1_FPCI_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.COMB.RSDECODE.UN1_FPCI_0_X\,
dataa => N_55,
datab => N_56,
datac => N_54);
GRLFPC20_V_STATE_0_SQMUXA_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111101111111")
port map (
combout => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
dataa => N_390,
datab => N_389,
datac => N_388);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC20.FPI.RST_0_G0_X\,
dataa => N_1,
datab => \GRLFPC20.R.MK.RST2\,
datac => \GRLFPC20.R.MK.RST\);
GRLFPC20_COMB_UN1_FPCI_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.COMB.UN1_FPCI_0_X\,
dataa => N_354,
datab => N_353,
datac => N_4);
GRLFPC20_R_A_RS1D_0_0_G4_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.R.A.RS1D_0_0_G4_1_X\,
dataa => N_49,
datab => N_48,
datac => N_52);
GRLFPC20_RS2_0_SQMUXA_0_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.RS2_0_SQMUXA_0_X\,
dataa => N_66,
datab => N_67,
datac => N_64);
GRLFPC20_COMB_FPDECODE_UN1_FPCI_7_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.UN1_FPCI_7_1_X\,
dataa => N_54,
datab => N_55,
datac => N_52);
GRLFPC20_R_A_MOV_RNO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000111")
port map (
combout => \GRLFPC20.R.A.MOV_0_0_G1_1_X\,
dataa => N_50,
datab => N_51,
datac => N_54);
GRLFPC20_N_1243_I_0_A2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.N_1243_I_0_A2_1_X\,
dataa => N_77,
datab => N_4,
datac => N_78);
GRLFPC20_R_MK_BUSY_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.R.MK.BUSY_0_0_G0_0_X\,
dataa => N_1,
datab => \GRLFPC20.R.MK.HOLDN1\,
datac => \GRLFPC20.R.MK.HOLDN2\);
GRLFPC20_R_MK_RST_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.COMB.V.MK.RST_1_0_G0_1_0_X\,
dataa => N_3,
datab => \GRLFPC20.R.MK.RST\,
datac => \GRLFPC20.R.MK.RST2\);
GRLFPC20_R_X_AFSR_RNISO6G: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.AFSR\,
datac => \GRLFPC20.R.X.LD\);
\GRLFPC20_WRDATA_X_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(14),
dataa => N_410,
datab => \GRLFPC20.WRDATA_0_X\(14),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(14),
dataa => N_410,
datab => \GRLFPC20.WRDATA_0_X\(46),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_RS1_1_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(2),
dataa => N_388,
datab => N_394,
datac => \GRLFPC20.COMB.RS1_1\(3));
\GRLFPC20_RS1_1_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(3),
dataa => N_388,
datab => N_395,
datac => \GRLFPC20.COMB.RS1_1\(4));
\GRLFPC20_RS2_1_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(3),
dataa => N_388,
datab => N_395,
datac => \GRLFPC20.COMB.RS2_1\(4));
\GRLFPC20_WRADDR_1_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => RFI2_WRADDRZ(2),
dataa => N_394,
datab => \GRLFPC20.WRADDR_0_SQMUXA_X\,
datac => \GRLFPC20.COMB.WRADDR_6_X\(3));
\GRLFPC20_WRADDR_1_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => RFI2_WRADDRZ(3),
dataa => N_395,
datab => \GRLFPC20.WRADDR_0_SQMUXA_X\,
datac => \GRLFPC20.COMB.WRADDR_6_X\(4));
\GRLFPC20_WRDATA_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(2),
dataa => N_398,
datab => \GRLFPC20.WRDATA_0_X\(2),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(11),
dataa => N_407,
datab => \GRLFPC20.WRDATA_0_X\(11),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(13),
dataa => N_409,
datab => \GRLFPC20.WRDATA_0_X\(13),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(17),
dataa => N_413,
datab => \GRLFPC20.WRDATA_0_X\(17),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(27),
dataa => N_423,
datab => \GRLFPC20.WRDATA_0_X\(27),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(29),
dataa => N_425,
datab => \GRLFPC20.WRDATA_0_X\(29),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(2),
dataa => N_398,
datab => \GRLFPC20.WRDATA_0_X\(34),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(11),
dataa => N_407,
datab => \GRLFPC20.WRDATA_0_X\(43),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(13),
dataa => N_409,
datab => \GRLFPC20.WRDATA_0_X\(45),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(17),
dataa => N_413,
datab => \GRLFPC20.WRDATA_0_X\(49),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(27),
dataa => N_423,
datab => \GRLFPC20.WRDATA_0_X\(59),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(29),
dataa => N_425,
datab => \GRLFPC20.WRDATA_0_X\(61),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRADDR_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => RFI2_WRADDRZ(0),
dataa => N_392,
datab => \GRLFPC20.WRADDR_0_SQMUXA_X\,
datac => \GRLFPC20.COMB.WRADDR_6_X\(1));
\GRLFPC20_WRADDR_1_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => RFI2_WRADDRZ(1),
dataa => N_393,
datab => \GRLFPC20.WRADDR_0_SQMUXA_X\,
datac => \GRLFPC20.COMB.WRADDR_6_X\(2));
\GRLFPC20_RS2_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(0),
dataa => N_388,
datab => N_392,
datac => \GRLFPC20.COMB.RS2_1\(1));
\GRLFPC20_WRDATA_X_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(21),
dataa => N_417,
datab => \GRLFPC20.WRDATA_0_X\(21),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(19),
dataa => N_415,
datab => \GRLFPC20.WRDATA_0_X\(19),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(18),
dataa => N_414,
datab => \GRLFPC20.WRDATA_0_X\(18),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(9),
dataa => N_405,
datab => \GRLFPC20.WRDATA_0_X\(9),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(6),
dataa => N_402,
datab => \GRLFPC20.WRDATA_0_X\(38),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(9),
dataa => N_405,
datab => \GRLFPC20.WRDATA_0_X\(41),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
GRLFPC20_COMB_ISFPOP2_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.COMB.ISFPOP2_1_X\,
dataa => N_338,
datab => \GRLFPC20.R.I.INST\(19),
datac => \GRLFPC20.COMB.UN1_R.I.V_0\);
\GRLFPC20_WRDATA_X_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(12),
dataa => N_408,
datab => \GRLFPC20.WRDATA_0_X\(12),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(15),
dataa => N_411,
datab => \GRLFPC20.WRDATA_0_X\(15),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(20),
dataa => N_416,
datab => \GRLFPC20.WRDATA_0_X\(20),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(23),
dataa => N_419,
datab => \GRLFPC20.WRDATA_0_X\(23),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(12),
dataa => N_408,
datab => \GRLFPC20.WRDATA_0_X\(44),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(15),
dataa => N_411,
datab => \GRLFPC20.WRDATA_0_X\(47),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(20),
dataa => N_416,
datab => \GRLFPC20.WRDATA_0_X\(52),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(23),
dataa => N_419,
datab => \GRLFPC20.WRDATA_0_X\(55),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_COMB_V_FSR_FCC_1_0_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC_1_0_X\(0),
dataa => N_406,
datab => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC20.R.I.CC\(0));
\GRLFPC20_COMB_V_FSR_FCC_1_0_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC_1_0_X\(1),
dataa => N_407,
datab => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC20.R.I.CC\(1));
\GRLFPC20_WRDATA_X_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(18),
dataa => N_414,
datab => \GRLFPC20.WRDATA_0_X\(50),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_RS2_1_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(2),
dataa => N_388,
datab => N_394,
datac => \GRLFPC20.COMB.RS2_1\(3));
\GRLFPC20_RS2_1_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD2ADDRZ(1),
dataa => N_388,
datab => N_393,
datac => \GRLFPC20.COMB.RS2_1\(2));
\GRLFPC20_WRDATA_X_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(8),
dataa => N_404,
datab => \GRLFPC20.WRDATA_0_X\(8),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(8),
dataa => N_404,
datab => \GRLFPC20.WRDATA_0_X\(40),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
GRLFPC20_V_FSR_NONSTD_0_SQMUXA_2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.AFSR\,
datac => \GRLFPC20.R.X.LD\);
\GRLFPC20_COMB_V_I_RES_6_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000010010")
port map (
combout => \GRLFPC20.COMB.V.I.RES_6_X\(63),
dataa => N_119,
datab => N_120,
datac => \GRLFPC20.FPI.OP2_X\(63));
\GRLFPC20_WRDATA_X_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(7),
dataa => N_403,
datab => \GRLFPC20.WRDATA_0_X\(7),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(10),
dataa => N_406,
datab => \GRLFPC20.WRDATA_0_X\(10),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(24),
dataa => N_420,
datab => \GRLFPC20.WRDATA_0_X\(24),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(31),
dataa => N_427,
datab => \GRLFPC20.WRDATA_0_X\(31),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(4),
dataa => N_400,
datab => \GRLFPC20.WRDATA_0_X\(36),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(7),
dataa => N_403,
datab => \GRLFPC20.WRDATA_0_X\(39),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(10),
dataa => N_406,
datab => \GRLFPC20.WRDATA_0_X\(42),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(24),
dataa => N_420,
datab => \GRLFPC20.WRDATA_0_X\(56),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(31),
dataa => N_427,
datab => \GRLFPC20.WRDATA_0_X\(63),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_R_X_SEQERR_RNIFJ4S_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101110101011")
port map (
combout => \GRLFPC20.UN1_FPCI_22_X\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.FPOP\,
datac => \GRLFPC20.R.X.SEQERR\(0));
\GRLFPC20_WRDATA_X_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(30),
dataa => N_426,
datab => \GRLFPC20.WRDATA_0_X\(62),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(1),
dataa => N_397,
datab => \GRLFPC20.WRDATA_0_X\(33),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(30),
dataa => N_426,
datab => \GRLFPC20.WRDATA_0_X\(30),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(28),
dataa => N_424,
datab => \GRLFPC20.WRDATA_0_X\(60),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(21),
dataa => N_417,
datab => \GRLFPC20.WRDATA_0_X\(53),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(28),
dataa => N_424,
datab => \GRLFPC20.WRDATA_0_X\(28),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(22),
dataa => N_418,
datab => \GRLFPC20.WRDATA_0_X\(22),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(19),
dataa => N_415,
datab => \GRLFPC20.WRDATA_0_X\(51),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(22),
dataa => N_418,
datab => \GRLFPC20.WRDATA_0_X\(54),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(0),
dataa => N_396,
datab => \GRLFPC20.WRDATA_0_X\(0),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(1),
dataa => N_397,
datab => \GRLFPC20.WRDATA_0_X\(1),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(5),
dataa => N_401,
datab => \GRLFPC20.WRDATA_0_X\(5),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_RS1_1_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(1),
dataa => N_388,
datab => N_393,
datac => \GRLFPC20.COMB.RS1_1\(2));
\GRLFPC20_WRDATA_X_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(26),
dataa => N_422,
datab => \GRLFPC20.WRDATA_0_X\(58),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(26),
dataa => N_422,
datab => \GRLFPC20.WRDATA_0_X\(26),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(25),
dataa => N_421,
datab => \GRLFPC20.WRDATA_0_X\(57),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(5),
dataa => N_401,
datab => \GRLFPC20.WRDATA_0_X\(37),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(0),
dataa => N_396,
datab => \GRLFPC20.WRDATA_0_X\(32),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(25),
dataa => N_421,
datab => \GRLFPC20.WRDATA_0_X\(25),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(4),
dataa => N_400,
datab => \GRLFPC20.WRDATA_0_X\(4),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_RS1_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => RFI2_RD1ADDRZ(0),
dataa => N_388,
datab => N_392,
datac => \GRLFPC20.COMB.RS1_1\(1));
\GRLFPC20_WRDATA_X_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(16),
dataa => N_412,
datab => \GRLFPC20.WRDATA_0_X\(48),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI1_WRDATAZ(3),
dataa => N_399,
datab => \GRLFPC20.WRDATA_0_X\(35),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(16),
dataa => N_412,
datab => \GRLFPC20.WRDATA_0_X\(16),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(6),
dataa => N_402,
datab => \GRLFPC20.WRDATA_0_X\(6),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
\GRLFPC20_WRDATA_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => RFI2_WRDATAZ(3),
dataa => N_399,
datab => \GRLFPC20.WRDATA_0_X\(3),
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\);
GRLFPC20_WREN2_1_SQMUXA_1_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.WREN2_1_SQMUXA_1_1_X\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.SEQERR\(0),
datac => \GRLFPC20.COMB.UN1_R.I.EXC\);
\GRLFPC20_COMB_V_FSR_CEXC_1_2_A_X_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110100011101")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(0),
dataa => N_396,
datab => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC20.R.I.EXC\(0));
\GRLFPC20_COMB_V_FSR_CEXC_1_2_A_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110100011101")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(1),
dataa => N_397,
datab => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC20.R.I.EXC\(1));
\GRLFPC20_COMB_V_FSR_CEXC_1_2_A_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110100011101")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(2),
dataa => N_398,
datab => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC20.R.I.EXC\(2));
\GRLFPC20_COMB_V_FSR_CEXC_1_2_A_X_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110100011101")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(3),
dataa => N_399,
datab => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC20.R.I.EXC\(3));
\GRLFPC20_COMB_V_FSR_CEXC_1_2_A_X_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110100011101")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(4),
dataa => N_400,
datab => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datac => \GRLFPC20.R.I.EXC\(4));
GRLFPC20_COMB_SEQERR_UN7_OP_0_A2_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010110000")
port map (
combout => \GRLFPC20.COMB.SEQERR.UN7_OP_0_A2_X\,
dataa => N_62,
datab => N_63,
datac => \GRLFPC20.COMB.RDD_1.M14_0_A2_1\);
GRLFPC20_V_STATE_1_SQMUXA_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC20.V.STATE_1_SQMUXA_1_X\,
dataa => N_424,
datab => N_1,
datac => \GRLFPC20.V.STATE_0_SQMUXA_1_X\);
GRLFPC20_COMB_FPDECODE_FPOP2_0_A2_RNISPI51: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.R.A.MOV_0_0_G1_0_X\,
dataa => N_74,
datab => N_73,
datac => \GRLFPC20.COMB.FPDECODE.FPOP2_0_A2\);
GRLFPC20_R_X_FPOP_RNIM15L: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
dataa => N_3,
datab => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datac => \GRLFPC20.R.X.FPOP\);
GRLFPC20_RS1V_0_SQMUXA_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000011100000")
port map (
combout => \GRLFPC20.RS1V_0_SQMUXA_1_X\,
dataa => \GRLFPC20.COMB.RSDECODE.RS1V2_0\,
datab => \GRLFPC20.COMB.FPDECODE.RDD5_0_A3\,
datac => \GRLFPC20.COMB.FPDECODE.FPOP2_0_A2\);
GRLFPC20_COMB_V_A_LD_1_0_O2_RNIV4FL1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\,
dataa => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_TZ\,
datab => \GRLFPC20.COMB.V.A.LD_1_0_O2\);
GRLFPC20_R_MK_BUSY2_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.R.MK.BUSY2_0_0_G0_X\,
dataa => N_1,
datab => \GRLFPC20.R.MK.BUSY\,
datac => \GRLFPC20.R.MK.BUSY2_0_0_G3\);
GRLFPC20_COMB_WREN2_11_IV_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110011101100")
port map (
combout => \GRLFPC20.COMB.WREN2_11_IV_1_X\,
dataa => N_344,
datab => \GRLFPC20.WREN2_1_SQMUXA_1\,
datac => \GRLFPC20.WREN2_2_SQMUXA_1\);
GRLFPC20_COMB_UN7_RS1V_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.COMB.UN7_RS1V_X\,
dataa => \GRLFPC20.COMB.RS1D_1_U\,
datab => \GRLFPC20.COMB.RS1_1\(0));
GRLFPC20_COMB_UN1_RS1V_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC20.COMB.UN1_RS1V_X\,
dataa => \GRLFPC20.COMB.RS1D_1_U\,
datab => \GRLFPC20.COMB.RS1_1\(0));
\GRLFPC20_COMB_V_A_RF1REN_1_1_X_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.COMB.V.A.RF1REN_1_1_X\(1),
dataa => \GRLFPC20.COMB.RS1V_1_IV\,
datab => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\);
GRLFPC20_RIN_MK_LDOP_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.RIN.MK.LDOP_X\,
dataa => N_3,
datab => \GRLFPC20.RS2_0_SQMUXA\,
datac => \GRLFPC20.R.A.AFSR_0_0_G1_1\);
\GRLFPC20_COMB_RF2REN_1_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.RF2REN_1_0_X\(2),
dataa => N_3,
datab => \GRLFPC20.R.A.RF2REN\(2),
datac => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I\);
\GRLFPC20_COMB_RF1REN_1_0_X_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.COMB.RF1REN_1_0_X\(2),
dataa => N_3,
datab => \GRLFPC20.R.A.RF1REN\(2),
datac => \GRLFPC20.COMB.V.A.RF1REN_1\(2));
GRLFPC20_COMB_WREN1_11_IV_1_X: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010110000")
port map (
combout => \GRLFPC20.COMB.WREN1_11_IV_1_X\,
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.COMB.WRADDR_6_X\(0),
datac => \GRLFPC20.COMB.WREN129\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_0_7__G0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010010000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_31_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31_S_0\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_S\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_27\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31_D\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_SCTRL_39_IV_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_1\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT_I_M\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN29_GRFPUSX_M_381\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV_0\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_A5_0_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_1__G0\,
dataa => N_52,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_1__G0_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_31_D_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31_D\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_15\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0\(75));
GRLFPC20_COMB_WREN1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011101000110000")
port map (
combout => RFI1_WRENZ,
dataa => N_3,
datab => N_391,
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\,
datad => \GRLFPC20.COMB.WREN1_11_IV\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_114__G0\,
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_114__G0_A\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_114__G0_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(114),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(114));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_1__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN14_CONDITIONAL\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4\);
\GRLFPC20_R_FSR_AEXC_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001100")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_0__G1\,
dataa => \GRLFPC20.R.FSR.AEXC\(0),
datab => \GRLFPC20.R.FSR.AEXC_1_0_0__G1_0\,
datac => \GRLFPC20.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(0));
\GRLFPC20_R_FSR_AEXC_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001100")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_2__G1\,
dataa => \GRLFPC20.R.FSR.AEXC\(2),
datab => \GRLFPC20.R.FSR.AEXC_1_0_2__G1_0\,
datac => \GRLFPC20.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_IV_I_0_0__G0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
datab => NN_1,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN29_GRFPUSX_M_381\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_IV_I_0_0__G0_0\);
\GRLFPC20_R_FSR_AEXC_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001100")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_3__G1\,
dataa => \GRLFPC20.R.FSR.AEXC\(3),
datab => \GRLFPC20.R.FSR.AEXC_1_0_3__G1_0\,
datac => \GRLFPC20.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(3));
\GRLFPC20_R_FSR_AEXC_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001100")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_4__G1\,
dataa => \GRLFPC20.R.FSR.AEXC\(4),
datab => \GRLFPC20.R.FSR.AEXC_1_0_4__G1_0\,
datac => \GRLFPC20.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(4));
\GRLFPC20_R_FSR_AEXC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010001100")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_1__G1\,
dataa => \GRLFPC20.R.FSR.AEXC\(1),
datab => \GRLFPC20.R.FSR.AEXC_1_0_1__G1_0\,
datac => \GRLFPC20.V.FSR.AEXC_2_SQMUXA\,
datad => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_15_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_15\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_15_D\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_6\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_30_D_0_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010010110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0_D_0\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_21\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111111101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(60),
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_319__G3_0_X2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(60));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(59),
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_318__G3_0_X2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4_A\(56),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4_A\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\);
GRLFPC20_COMB_WREN2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011000000")
port map (
combout => RFI2_WRENZ,
dataa => N_3,
datab => N_391,
datac => \GRLFPC20.WRADDR_0_SQMUXA_X\,
datad => \GRLFPC20.COMB.WREN2_11_IV\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_SCTRL_39_IV_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(0),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.FPI.OP2_X\(63),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_0\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101011001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_IV_I_0_0__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
datab => \GRLFPC20.FPI.OP1_X\(63),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_AREGSIGN_SEL_30\);
GRLFPC20_COMB_WREN1_11_IV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111011100")
port map (
combout => \GRLFPC20.COMB.WREN1_11_IV\,
dataa => N_344,
datab => \GRLFPC20.WREN1_1_SQMUXA\,
datac => \GRLFPC20.WREN2_2_SQMUXA_1\,
datad => \GRLFPC20.COMB.WREN1_11_IV_1_X\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN20_STKOUT_RNIOBJES: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_S\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_15_D_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_15_D\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_14\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_3\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_30_D_0_D_0_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0_D_0\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0_D\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_18\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(58),
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.CO0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_27_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_27\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN14_CONDITIONAL\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_A5_0_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1\);
\GRLFPC20_R_FSR_AEXC_RNO_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011111010")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_4__G1_0\,
dataa => N_405,
datab => N_365,
datac => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC20.V.FSR.AEXC_1_SQMUXA\);
\GRLFPC20_R_FSR_AEXC_RNO_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011111010")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_2__G1_0\,
dataa => N_403,
datab => N_363,
datac => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC20.V.FSR.AEXC_1_SQMUXA\);
\GRLFPC20_R_FSR_AEXC_RNO_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011111010")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_1__G1_0\,
dataa => N_402,
datab => N_362,
datac => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC20.V.FSR.AEXC_1_SQMUXA\);
\GRLFPC20_R_FSR_AEXC_RNO_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011111010")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_3__G1_0\,
dataa => N_404,
datab => N_364,
datac => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC20.V.FSR.AEXC_1_SQMUXA\);
\GRLFPC20_R_FSR_AEXC_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011111010")
port map (
combout => \GRLFPC20.R.FSR.AEXC_1_0_0__G1_0\,
dataa => N_401,
datab => N_361,
datac => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datad => \GRLFPC20.V.FSR.AEXC_1_SQMUXA\);
\GRLFPC20_R_FSR_AEXC_RNO_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(0),
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.R.FSR.AEXC\(0),
datac => \GRLFPC20.R.I.EXC\(0),
datad => \GRLFPC20.R.I.V_EN_1\);
\GRLFPC20_R_FSR_AEXC_RNO_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(2),
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.R.FSR.AEXC\(2),
datac => \GRLFPC20.R.I.EXC\(2),
datad => \GRLFPC20.R.I.V_EN_1\);
\GRLFPC20_R_FSR_AEXC_RNO_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(3),
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.R.FSR.AEXC\(3),
datac => \GRLFPC20.R.I.EXC\(3),
datad => \GRLFPC20.R.I.V_EN_1\);
\GRLFPC20_R_FSR_AEXC_RNO_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(4),
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.R.FSR.AEXC\(4),
datac => \GRLFPC20.R.I.EXC\(4),
datad => \GRLFPC20.R.I.V_EN_1\);
\GRLFPC20_R_FSR_AEXC_RNO_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.COMB.V.FSR.AEXC_7_I_M\(1),
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.R.FSR.AEXC\(1),
datac => \GRLFPC20.R.I.EXC\(1),
datad => \GRLFPC20.R.I.V_EN_1\);
GRLFPC20_COMB_WREN2_11_IV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011110000")
port map (
combout => \GRLFPC20.COMB.WREN2_11_IV\,
dataa => \GRLFPC20.COMB.RDD_2\,
datab => \GRLFPC20.COMB.WRADDR_6_X\(0),
datac => \GRLFPC20.COMB.WREN2_11_IV_1_X\,
datad => \GRLFPC20.COMB.WREN129\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_SCTRL_39_IV_0_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_0\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_0_A\(12),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_SCTRL_39_IV_0_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_0_A\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.UN4_TEMP\,
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_E\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_18_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101101000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_18\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_RNI2FG5C_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_318__G3_0_X2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_0_A2\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_261__G5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN2_MIXOIN_25_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110011101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19_U\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_316_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_316__G3_0_X2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_9\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_BNC4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_259__G5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_3_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_3\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_RNI0H7CE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_319__G3_0_X2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_ANC3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.CO0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN30_CONDITIONAL_0_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(9));
GRLFPC20_R_I_V_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.R.I.V_1_0_G0_0\,
dataa => \GRLFPC20.COMB.UN1_R.I.EXC\,
datab => \GRLFPC20.COMB.ANNULRES_1_IV_454\,
datac => \GRLFPC20.R.I.V_1_0_G0_0_1\,
datad => \GRLFPC20.R.I.V_EN_1\);
GRLFPC20_V_FSR_CEXC_3_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\,
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\,
datac => \GRLFPC20.COMB.V.STATE14\,
datad => \GRLFPC20.R.I.V_EN_1\);
GRLFPC20_R_I_EXEC_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.R.I.EXEC_0_0_G1_0_549_I\,
dataa => \GRLFPC20.R.I.EXEC_0_0_G1_0_I_0_0\,
datab => \GRLFPC20.R.I.EXEC_0_0_G1_0_I_A8_0\,
datac => \GRLFPC20.COMB.ANNULRES_1_IV_454\,
datad => \GRLFPC20.R.I.V_EN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_WQSCTRL_RNILHL93_0_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT_0\(1));
GRLFPC20_V_FSR_AEXC_2_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.V.FSR.AEXC_2_SQMUXA\,
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\,
datac => \GRLFPC20.COMB.V.FSR.FCC10\,
datad => \GRLFPC20.COMB.WREN129\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_XZBREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_E\);
GRLFPC20_V_FSR_AEXC_1_SQMUXA_0_RNIL956: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111101")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M3\,
dataa => \GRLFPC20.V.FSR.AEXC_1_SQMUXA_0\,
datab => \GRLFPC20.COMB.V.STATE14\,
datac => \GRLFPC20.COMB.V.FSR.FCC10\,
datad => \GRLFPC20.V.FSR.CEXC_3_SQMUXA\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0_A2\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_WQSCTRL_RNIENRC2_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN29_GRFPUSX_M_381\,
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN2_AREGSIGN_SEL_30: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_AREGSIGN_SEL_30\,
dataa => NN_1,
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_E\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_XZAREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_COMB_RF1REN_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI1_REN2Z,
dataa => N_390,
datab => N_389,
datac => N_388,
datad => \GRLFPC20.COMB.RF1REN_1_0_X\(2));
\GRLFPC20_COMB_V_FSR_FCC_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110011100100")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC_1\(1),
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.COMB.V.FSR.FCC_1_0_X\(1),
datac => \GRLFPC20.COMB.V.FSR.FCC_1_1_X\(1),
datad => \GRLFPC20.COMB.V.FSR.FCC10\);
\GRLFPC20_COMB_V_FSR_FCC_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110011100100")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC_1\(0),
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.COMB.V.FSR.FCC_1_0_X\(0),
datac => \GRLFPC20.COMB.V.FSR.FCC_1_1_X\(0),
datad => \GRLFPC20.COMB.V.FSR.FCC10\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_23_1_CO0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.CO0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.CO0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.SUM_0_A2\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_51\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_53\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_52\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_54\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_RNI2FG5C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_0_A2\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_261__G5\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN36_STKGEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110100000010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_SCTRL_39_IV_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT_I_M\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT_I_M_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
GRLFPC20_R_MK_BUSY_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC20.R.MK.BUSY_0_0_G0\,
dataa => \GRLFPC20.R.MK.BUSY_0_0_G0_0_X\,
datab => \GRLFPC20.FPI.LDOP_2\,
datac => \GRLFPC20.R.MK.BUSY2_0_0_G3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP\);
GRLFPC20_R_MK_RST_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.COMB.V.MK.RST_1_0_G0\,
dataa => \GRLFPC20.COMB.V.MK.RST_1_0_G0_1_0_X\,
datab => CPO_HOLDNZ,
datac => \GRLFPC20.R.MK.BUSY2_0_0_G3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_8_1_SUM_0_A2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0_A2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_9\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_BNC4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_259__G5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_23_1_SUM_0_A2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.SUM_0_A2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.CO0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_258_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_258__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.CO0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_0_A2\(56));
GRLFPC20_V_FSR_AEXC_1_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010001000")
port map (
combout => \GRLFPC20.V.FSR.AEXC_1_SQMUXA\,
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\,
datac => \GRLFPC20.COMB.ISFPOP2_1_X\,
datad => \GRLFPC20.COMB.V.FSR.FCC10_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3_RNIK5TVA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011111101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_14_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010011010010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_14\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_12\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_9\(75));
\GRLFPC20_COMB_RF2REN_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI2_REN2Z,
dataa => N_390,
datab => N_389,
datac => N_388,
datad => \GRLFPC20.COMB.RF2REN_1_0_X\(2));
\GRLFPC20_COMB_RF1REN_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI1_REN1Z,
dataa => N_390,
datab => N_389,
datac => N_388,
datad => \GRLFPC20.COMB.RF1REN_1_0\(1));
\GRLFPC20_COMB_RF2REN_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111110110000")
port map (
combout => RFI2_REN1Z,
dataa => N_390,
datab => N_389,
datac => N_388,
datad => \GRLFPC20.COMB.RF2REN_1_0\(1));
GRLFPC20_COMB_V_FSR_FCC10_1_RNI2I2J: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000011010000")
port map (
combout => \GRLFPC20.R.I.V_EN_1\,
dataa => \GRLFPC20.R.X.LD\,
datab => \GRLFPC20.COMB.ISFPOP2_1_X\,
datac => \GRLFPC20.COMB.V.FSR.FCC10_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN30_CONDITIONAL_0_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000110010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN12_STKOUT_RNIUR8UA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_STKOUT\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0\,
dataa => N_53,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0\);
\GRLFPC20_COMB_V_A_RF1REN_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010000000000")
port map (
combout => \GRLFPC20.COMB.V.A.RF1REN_1\(2),
dataa => N_43,
datab => \GRLFPC20.RS2_0_SQMUXA\,
datac => \GRLFPC20.COMB.RS2D_1_IV\,
datad => \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2\);
GRLFPC20_COMB_WREN129: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.COMB.WREN129\,
dataa => \GRLFPC20.R.X.LD\,
datab => \GRLFPC20.COMB.ISFPOP2_1_X\,
datac => \GRLFPC20.COMB.V.FSR.FCC10_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_BUSYMULXFF_UN2_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_8_1_SUM_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_ANC3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.CO0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_PCTRL_NEW_43_1_RNIJ1GT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110011101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_8_RNIIQ021: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010111110001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL_1_0\(67),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(173),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(57));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN20_STKOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101101011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN20_STKOUT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN2_MIXOIN_19_U_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_19_U\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_CI_114_1_CO0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.CO0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN38_PCTRL_NEW_I_0_G0\,
dataa => \GRLFPC20.FPI.LDOP_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20\,
datac => \GRLFPC20.RIN.MK.LDOP_X\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_6_0_67__G0_E_I\,
dataa => N_3,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datac => \GRLFPC20.FPI.LDOP_2\,
datad => \GRLFPC20.R.A.FPOP_0_0_G1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_RESULT_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT_0\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\);
\GRLFPC20_COMB_RF2REN_1_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010001000100")
port map (
combout => \GRLFPC20.COMB.RF2REN_1_0\(1),
dataa => N_3,
datab => \GRLFPC20.R.A.RF2REN\(1),
datac => \GRLFPC20.COMB.UN7_RS1V_X\,
datad => \GRLFPC20.COMB.V.A.RF1REN_1_1_X\(1));
\GRLFPC20_COMB_RF1REN_1_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010001000100")
port map (
combout => \GRLFPC20.COMB.RF1REN_1_0\(1),
dataa => N_3,
datab => \GRLFPC20.R.A.RF1REN\(1),
datac => \GRLFPC20.COMB.UN1_RS1V_X\,
datad => \GRLFPC20.COMB.V.A.RF1REN_1_1_X\(1));
GRLFPC20_COMB_V_FSR_FCC10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC10\,
dataa => \GRLFPC20.COMB.ISFPOP2_1_X\,
datab => \GRLFPC20.COMB.UN1_R.I.V\,
datac => \GRLFPC20.COMB.V.STATE\,
datad => \GRLFPC20.R.STATE_0_0_0__G3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_1\,
dataa => N_54,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_A5_0_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_A\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0_0_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_52: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_52\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_11\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_35\);
\GRLFPC20_R_A_RF1REN_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110000000000")
port map (
combout => \GRLFPC20.COMB.V.A.RF1REN_1_670_I\,
dataa => \GRLFPC20.COMB.RS1D_1_U\,
datab => \GRLFPC20.COMB.RS1V_1_IV\,
datac => \GRLFPC20.COMB.V.A.RF1REN_1_670_I_M4\,
datad => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\);
\GRLFPC20_R_A_RF2REN_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000000")
port map (
combout => \GRLFPC20.COMB.V.A.RF2REN_1_734_I\,
dataa => \GRLFPC20.COMB.RS1D_1_U\,
datab => \GRLFPC20.COMB.RS1V_1_IV\,
datac => \GRLFPC20.COMB.V.A.RF1REN_1_670_I_M4\,
datad => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\);
\GRLFPC20_R_STATE_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110000000000")
port map (
combout => \GRLFPC20.R.STATE_0_0_0__G1\,
dataa => N_5,
datab => \GRLFPC20.V.STATE_1_SQMUXA_1_X\,
datac => CPO_EXCZ,
datad => \GRLFPC20.R.STATE_0_0_0__G3\);
GRLFPC20_COMB_V_FSR_FCC10_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.COMB.V.FSR.FCC10_1\,
dataa => \GRLFPC20.COMB.UN1_R.I.V\,
datab => \GRLFPC20.COMB.V.STATE\,
datac => \GRLFPC20.R.STATE_0_0_0__G3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_BUSYMULXFF_UN2_TEMP_1_RNIQG4O3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_10_RNI571R5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000011110110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_261__G5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.ANC1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_CI_114_1_SUM_0_A2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100010000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_0_A2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_TEMP_RNIVRVM5_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN22_NOTPROP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM1_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN19_GEN\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_3_RNIH2UH4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_259__G5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_9_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_9\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\);
GRLFPC20_FPI_START: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.FPI.START\,
dataa => N_3,
datab => \GRLFPC20.RS2_0_SQMUXA\,
datac => \GRLFPC20.FPI.LDOP_2\,
datad => \GRLFPC20.R.A.AFSR_0_0_G1_1\);
GRLFPC20_COMB_RS2D_1_IV_RNIR8PB2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000000000")
port map (
combout => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I\,
dataa => N_43,
datab => \GRLFPC20.RS2_0_SQMUXA\,
datac => \GRLFPC20.COMB.RS2D_1_IV\,
datad => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\);
\GRLFPC20_R_STATE_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010000000")
port map (
combout => \GRLFPC20.R.STATE_0_0_1__G1\,
dataa => N_5,
datab => \GRLFPC20.V.STATE_1_SQMUXA_1_X\,
datac => CPO_EXCZ,
datad => \GRLFPC20.COMB.V.STATE\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_53_SI_118_1_CO0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110100011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.CO0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_SUM2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.CO0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3_RNIPCSJ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100010000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_0_A2\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\(56));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_BUSYMULXFF_UN2_TEMP_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(70),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_65__G3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN4_STKOUT_RNIPBJK7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0_A3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN4_STKOUT\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOINSTANDNOEXC_41_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_PCTRL_NEW_43_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN27_STKGEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001011001101001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_V\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN27_STKGEN_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN27_STKGEN_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_0\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_10_RNI571R5_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001011001101001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.ANC1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\(56));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSAMPLEDWAIT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\);
\GRLFPC20_R_STATE_RNIES063_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011110000")
port map (
combout => \GRLFPC20.R.STATE_0_0_0__G3\,
dataa => \GRLFPC20.R.STATE\(0),
datab => \GRLFPC20.UN1_FPCI_2\,
datac => \GRLFPC20.R.STATE_0_0_0__G3_0\,
datad => \GRLFPC20.R.FSR.FTT_1_0_2__G2_490\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_53_SI_118_1_SUM_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001011010010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.SUM\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_SUM2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.CO0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(57),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN19_GEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN19_GEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM1_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C1_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_RNI486R4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_V\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_3_RNI014I2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_BNC4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C2\);
\GRLFPC20_R_I_EXC_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000010")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_2__G0\,
dataa => \GRLFPC20.R.I.EXC\(2),
datab => \GRLFPC20.COMB.UN2_HOLDN\,
datac => \GRLFPC20.COMB.UN19_IUEXEC\,
datad => \GRLFPC20.R.I.EXC_2_0_2__G3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0_A5_0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529_A3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_35: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_35\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(45),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_35_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_35_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100011111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_35_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(40),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_4\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_1_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0\,
dataa => N_49,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0\);
GRLFPC20_R_A_AFSR_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC20.R.A.AFSR_0_0_G1\,
dataa => N_66,
datab => \GRLFPC20.R.A.AFSR_0_0_G1_1_0\,
datac => \GRLFPC20.COMB.FPDECODE.FPOP8_I_O3_X\,
datad => \GRLFPC20.R.A.AFSR_0_0_G1_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_2__G0\,
dataa => N_50,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_2__G0_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101111111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_65__G0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529_A3\);
GRLFPC20_R_A_AFQ_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.R.A.AFQ_0_0_G1\,
dataa => \GRLFPC20.N_1243_I_0_A2_1_X\,
datab => \GRLFPC20.R.A.AFQ_0_0_G1_0\,
datac => CPO_EXCZ,
datad => \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2_RNIANRT1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_RNITGSH2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(12),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(13),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(40),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(42),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(44),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(48),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(50),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(49),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(51),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(11),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(14),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(17),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(19),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(20),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(22),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(24),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(25),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(26),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(28),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(30),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(33),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(37),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(38),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(39),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(41),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(18),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(21),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(23),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(27),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(36),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(47),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(52),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(45),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(15),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(15));
GRLFPC20_R_I_V_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC20.R.I.V_1_0_G3\,
dataa => \GRLFPC20.COMB.UN1_R.I.EXC\,
datab => \GRLFPC20.COMB.V.I.V_1_F1\,
datac => \GRLFPC20.COMB.ANNULRES_1_IV_454\);
GRLFPC20_COMB_RS2D_1_IV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011000000")
port map (
combout => \GRLFPC20.COMB.RS2D_1_IV\,
dataa => \GRLFPC20.COMB.V.A.RF1REN_1_0_650_A2_3_X\,
datab => \GRLFPC20.MOV_7_SQMUXA\,
datac => \GRLFPC20.R.A.RS1D_0_0_G4\,
datad => \GRLFPC20.UN1_MOV_1_SQMUXA\);
GRLFPC20_COMB_RS1V_1_IV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC20.COMB.RS1V_1_IV\,
dataa => \GRLFPC20.RS1V_0_SQMUXA\,
datab => \GRLFPC20.COMB.RSDECODE.RS1V_X\,
datac => \GRLFPC20.COMB.V.A.RF1REN_1_0_650_A2_3_X\,
datad => \GRLFPC20.UN1_RS1V_0_SQMUXA\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(55));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_RNI7N992: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN12_STKOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000111111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN12_STKOUT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0_A3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_STKGEN\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN2_MIXOIN_9_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_9\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0_A3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(43),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(53),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(46),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(54),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(54));
GRLFPC20_COMB_V_A_AFSR_1_5_0_O2_RNIVSQN1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.R.A.FPOP_0_0_G1\,
dataa => \GRLFPC20.N_1243_I_0_A2_1_X\,
datab => \GRLFPC20.RS2_0_SQMUXA\,
datac => CPO_EXCZ,
datad => \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2\);
\GRLFPC20_R_A_RDD_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC20.R.A.RDD_0_0_0__G1_0\,
dataa => N_62,
datab => N_63,
datac => \GRLFPC20.COMB.RDD_1.M14_0_A2_1\,
datad => \GRLFPC20.R.A.RDD_0_0_0__G2\);
GRLFPC20_V_FSR_FTT_1_SQMUXA_0_RNIPMDG2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110011001100")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_0__G0_I_O4_I\,
dataa => N_1,
datab => N_3,
datac => \GRLFPC20.UN1_FPCI_13\,
datad => \GRLFPC20.R.FSR.FTT_1_0_2__G2_490\);
GRLFPC20_COMB_V_STATE14_RNIBI0N1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.COMB.V.STATE\,
dataa => \GRLFPC20.R.STATE\(1),
datab => \GRLFPC20.UN1_FPCI_2\,
datac => \GRLFPC20.COMB.V.STATE14\,
datad => \GRLFPC20.COMB.UN1_R.I.EXC\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNISM4Q1_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_65__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529_A3\);
\GRLFPC20_R_I_EXC_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000000010")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_0__G0\,
dataa => \GRLFPC20.R.I.EXC\(0),
datab => \GRLFPC20.COMB.UN2_HOLDN\,
datac => \GRLFPC20.COMB.UN19_IUEXEC\,
datad => \GRLFPC20.R.I.EXC_2_0_0__G4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(35),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(29),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_2__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN14_CONDITIONAL\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_54: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_40\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_41\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_50\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_53: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_53\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_38\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_39\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_47\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000010010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_5\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_9_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_9_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_9_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_2\);
GRLFPC20_R_I_V_RNO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111101")
port map (
combout => \GRLFPC20.R.I.V_1_0_G0_0_1\,
dataa => N_1,
datab => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_A6_1_0\,
datac => \GRLFPC20.COMB.V.STATE14\,
datad => \GRLFPC20.G_884\);
GRLFPC20_COMB_V_STATE14_RNIKJ7T: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC20.R.STATE_0_0_0__G3_0\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.SEQERR\(0),
datac => \GRLFPC20.COMB.V.STATE14\,
datad => \GRLFPC20.COMB.UN1_R.I.EXC\);
\GRLFPC20_R_I_EXC_RNO_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_2__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
datac => \GRLFPC20.COMB.UN2_HOLDN\,
datad => \GRLFPC20.R.I.EXC_2_0_0__G4\);
\GRLFPC20_R_A_SEQERR_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC20.R.A.SEQERR_0_0_0__G1\,
dataa => \GRLFPC20.N_1243_I_0_A2_1_X\,
datab => CPO_EXCZ,
datac => \GRLFPC20.R.A.SEQERR_0_0_0__G3\,
datad => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\);
\GRLFPC20_R_A_RDD_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.R.A.RDD_0_0_0__G2\,
dataa => N_56,
datab => N_52,
datac => \GRLFPC20.COMB.RDD_1.M14_0_O2\,
datad => \GRLFPC20.R.A.MOV_0_0_G1_0_X\);
\GRLFPC20_R_FSR_FTT_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_2__G2\,
dataa => N_1,
datab => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_A6_1_0\,
datac => \GRLFPC20.COMB.V.STATE14\,
datad => \GRLFPC20.COMB.UN1_R.I.EXC\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(7));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN19_GEN_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C1_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(5),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011110010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(9),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(45));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000001010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(57),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_0_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_0_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRONEMORE\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN7_SHDVAR\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(57),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(15));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2_RNIANRT1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_SUM2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_54_SI_61_1_CO0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.CO0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_AXB0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_CI_58_2_ANC1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_58_2.ANC1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_1_RNIH1QV1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100010000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.SI_1_0_A2\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\(0));
GRLFPC20_COMB_RS1D_1_U: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011000000")
port map (
combout => \GRLFPC20.COMB.RS1D_1_U\,
dataa => \GRLFPC20.RS1D_CNST_0_A2_1_X\,
datab => \GRLFPC20.MOV_7_SQMUXA\,
datac => \GRLFPC20.R.A.RS1D_0_0_G4\,
datad => \GRLFPC20.RS1D_CNST_0_A2_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN19_GEN_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001000101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_0\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_1_RNIIO8B2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN16_NOTPROP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_0\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(7),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(55));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_GEN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.GEN_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM_I\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN13_GEN_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2_RNIDECL1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(54));
GRLFPC20_COMB_V_A_AFSR_1_5_0_O2_RNICIAC1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001000000000")
port map (
combout => \GRLFPC20.R.A.AFSR_0_0_G1_1\,
dataa => \GRLFPC20.N_1243_I_0_A2_1_X\,
datab => \GRLFPC20.R.STATE\(0),
datac => \GRLFPC20.R.STATE\(1),
datad => \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_STARTSHFT_UN3_NOTRESETORUNIMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000111110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529_A3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529_A3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001011010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_51: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_51\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_45\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_44\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_50: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_28\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_42\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_47: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_47\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_16\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_17\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_14\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_15\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_8\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(11));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(14),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(12));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101101111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_10_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_10_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111101101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(9),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_2\);
GRLFPC20_UN1_MOV_1_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111101000000")
port map (
combout => \GRLFPC20.UN1_MOV_1_SQMUXA\,
dataa => N_56,
datab => \GRLFPC20.COMB.FPDECODE.RDD3_TZ\,
datac => \GRLFPC20.COMB.FPDECODE.FPOP2_0_A2\,
datad => \GRLFPC20.UN1_MOV_1_SQMUXA_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_374_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110011111000011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_374__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_374__G0_0_A\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_374_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000101000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_374__G0_0_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_54_SI_61_1_SUM_0_A2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.SUM_0_A2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_AXB0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN18_STKGEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001011010010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN18_STKGEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM_I\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_OPREXC_RNIUUGR1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_1\(77),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXC\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN13_EXMIPTRLSBS_M\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\);
GRLFPC20_COMB_UN1_R_I_EXC_RNIH7PC3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110011111")
port map (
combout => \GRLFPC20.COMB.ANNULRES_1_IV_454\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.COMB.ANNULRES_1_IV_454_A\,
datac => \GRLFPC20.ANNULRES_1_SQMUXA\,
datad => \GRLFPC20.COMB.UN1_R.I.EXC\);
\GRLFPC20_R_X_SEQERR_RNIPUP91_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100000101")
port map (
combout => \GRLFPC20.COMB.ANNULRES_1_IV_454_A\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.I.EXEC\,
datac => \GRLFPC20.R.X.SEQERR\(0),
datad => \GRLFPC20.R.X.FPOP\);
GRLFPC20_R_A_LD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.R.A.LD_0_0_G1\,
dataa => \GRLFPC20.N_1243_I_0_A2_1_X\,
datab => \GRLFPC20.COMB.SEQERR.UN7_OP_0_A2_X\,
datac => CPO_EXCZ,
datad => \GRLFPC20.COMB.V.A.LD_1_0_O2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_ENTRYPOINT_2_RNI6OD31: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529_A3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_ENTRYPOINT\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_5_A\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_5_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_30_D_0_D_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_D_0_D\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_25\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_S\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN14_CONDITIONAL\);
GRLFPC20_UN1_RS1V_0_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110000000")
port map (
combout => \GRLFPC20.UN1_RS1V_0_SQMUXA\,
dataa => N_62,
datab => N_64,
datac => \GRLFPC20.COMB.FPDECODE.FPOP3_0\,
datad => \GRLFPC20.RS1V_0_SQMUXA_1_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(12),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(13),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(40),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(42),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(44),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(48),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(50),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(27),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(49),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(51),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(56),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(11),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(14),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(17),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(19),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(20),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(22),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(24),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(25),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(26),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(28),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(30),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(33),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(37),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(38),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(39),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(41),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(52),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(18),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(21),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(23),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(36),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(47),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(45),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_141_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(141),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(141),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(141));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(15),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(15));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_10_RNILR0C1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.CO0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7356\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_5_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(116),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(55));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_1_RNITIDS5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100110010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(43),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(53),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(46),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(54),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(54));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_RNIKLT32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110010001100")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_0__G4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STATUS\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN3_INEXACT\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT\);
GRLFPC20_COMB_V_A_AFSR_1_5_0_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100000010")
port map (
combout => \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2\,
dataa => \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2_1\,
datab => \GRLFPC20.COMB.FPDECODE.ST_0_A2\,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.COMB.V.A.LD_1_0_O2\);
GRLFPC20_COMB_V_I_EXEC_5_IV_RNIUB4S: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011011111")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_2__G2_490\,
dataa => \GRLFPC20.R.I.V\,
datab => \GRLFPC20.COMB.UN1_MEXC_1\,
datac => \GRLFPC20.COMB.V.I.EXEC_5_IV\,
datad => \GRLFPC20.COMB.UN1_R.I.EXC\);
GRLFPC20_COMB_UN1_R_I_EXC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.COMB.UN1_R.I.EXC\,
dataa => \GRLFPC20.R.I.V\,
datab => \GRLFPC20.R.I.EXC\(5),
datac => \GRLFPC20.COMB.UN1_MEXC_1\,
datad => \GRLFPC20.COMB.V.I.EXEC_5_IV\);
GRLFPC20_COMB_V_I_EXEC_5_IV_RNIUN111: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M2\,
dataa => \GRLFPC20.V.STATE_0_SQMUXA_1_X\,
datab => \GRLFPC20.R.I.V\,
datac => \GRLFPC20.COMB.UN1_MEXC_1\,
datad => \GRLFPC20.COMB.V.I.EXEC_5_IV\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(35),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(29),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_SCTRL_39_IV_RNO_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT_I_M_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT\,
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_45: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_45\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_32\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_44: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_35\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_30\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_42: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_57\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_27\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_41: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_41\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_31\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_25\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_40: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_40\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_43\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_22\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_39: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_39\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_37\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_21\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_38: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_38\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_38\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_18\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110110110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(7),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(8));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOINSTANDNOEXC_41_2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTNULLEXC\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN13_GEN_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100010101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN13_GEN_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_2\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM0\);
GRLFPC20_RS1D_CNST_0_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010000000")
port map (
combout => \GRLFPC20.RS1D_CNST_0_A2_0\,
dataa => N_73,
datab => \GRLFPC20.RS1D_CNST_0_A2_0_A\,
datac => \GRLFPC20.RS1D_CNST_0_A2_2_X\,
datad => \GRLFPC20.COMB.FPDECODE.RDD5_0_A3\);
GRLFPC20_RS1D_CNST_0_A2_0_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000001100")
port map (
combout => \GRLFPC20.RS1D_CNST_0_A2_0_A\,
dataa => N_62,
datab => N_66,
datac => N_63,
datad => N_73);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_WAITMULXFF_NOTSAMPLEDWAIT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTNULLEXC\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.UN2_TEMP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS\(0));
GRLFPC20_COMB_V_I_EXEC_5_IV_RNINBKI: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.COMB.UN1_R.I.V\,
dataa => \GRLFPC20.R.I.V\,
datab => \GRLFPC20.COMB.UN1_MEXC_1\,
datac => \GRLFPC20.COMB.V.I.EXEC_5_IV\);
GRLFPC20_COMB_FPDECODE_ST3_1_RNI0EBA1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000001010001")
port map (
combout => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_TZ\,
dataa => \GRLFPC20.RS2_0_SQMUXA\,
datab => \GRLFPC20.COMB.FPDECODE.ST3_1\,
datac => \GRLFPC20.COMB.FPDECODE.FPOP8_I_O3_X\,
datad => \GRLFPC20.COMB.SEQERR.UN7_OP_0_A2_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI16741_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_C0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_RNI9HRN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_C0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI2TFQ_0_368_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_C0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_V\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(11));
GRLFPC20_COMB_RDD_1_M14_0_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111001101010000")
port map (
combout => \GRLFPC20.COMB.RDD_1.M14_0_O2\,
dataa => N_53,
datab => N_55,
datac => \GRLFPC20.COMB.RDD_1.M14_0_A2_0_0\,
datad => \GRLFPC20.COMB.RDD_1.M14_0_A2_0_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(5),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(9),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_14_141_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110000001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(141),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(143),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_171_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(171),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLCREGXZ.UN1_INFORCREGDB\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(171),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(7),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_NOTSRRES_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSRRES\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRONEMORE\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(54),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIGAOS4_370_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(370),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_2_I_O3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_10_RNIEA5N1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_10_RNIEA5N1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_ANC3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_BUSYMULXFF_UN2_TEMP_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.BUSYMULXFF.UN2_TEMP_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTNULLEXC\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_OPREXC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111101111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXC\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010000000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_A\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_4_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD11\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M5\);
GRLFPC20_COMB_V_A_LD_1_0_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011111110")
port map (
combout => \GRLFPC20.COMB.V.A.LD_1_0_O2\,
dataa => \GRLFPC20.COMB.RSDECODE.RS1V_X\,
datab => \GRLFPC20.COMB.LOCKGEN.LOCKI_I_0_0_A2_0\,
datac => \GRLFPC20.COMB.V.A.LD_1_0_A2_0\,
datad => \GRLFPC20.COMB.LOCKGEN.DEPCHECK\);
GRLFPC20_ANNULFPU_0_SQMUXA_1_X_RNI8NJG1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC20.R.MK.BUSY2_0_0_G3\,
dataa => \GRLFPC20.ANNULFPU_0_SQMUXA_1_X\,
datab => \GRLFPC20.ANNULFPU_0_SQMUXA_2_X\,
datac => \GRLFPC20.R.MK.BUSY2_0_0_G3_A\,
datad => \GRLFPC20.COMB.UN1_R.I.EXC\);
GRLFPC20_ANNULFPU_0_SQMUXA_X_RNIACM31: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100111")
port map (
combout => \GRLFPC20.R.MK.BUSY2_0_0_G3_A\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.FPOP\,
datac => \GRLFPC20.R.X.SEQERR\(0),
datad => \GRLFPC20.ANNULFPU_0_SQMUXA_X\);
GRLFPC20_COMB_V_STATE14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.COMB.V.STATE14\,
dataa => \GRLFPC20.R.I.V\,
datab => \GRLFPC20.COMB.UN1_MEXC_1\,
datac => \GRLFPC20.COMB.V.I.EXEC_5_IV\);
\GRLFPC20_R_A_SEQERR_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101011001100")
port map (
combout => \GRLFPC20.R.A.SEQERR_0_0_0__G3\,
dataa => \GRLFPC20.RS2_0_SQMUXA\,
datab => \GRLFPC20.R.A.AFQ_0_0_G1_0\,
datac => \GRLFPC20.COMB.SEQERR.UN7_OP_0_A2_X\,
datad => \GRLFPC20.COMB.QNE2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_32\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(46),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(18));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_30: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(23),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(17));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_29: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(26),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(21));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_28: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(24),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(16));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(47),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(34));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_25: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(28));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_22: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(56),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(48));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_21: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_21\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(54),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(53));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_18\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(39),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(33));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_17\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(52),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(30));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_16\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(44),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(20));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_15\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(51),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(41));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZZERO_1_14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010000100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZZERO_1_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(25),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(15));
GRLFPC20_R_I_EXEC_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010000000")
port map (
combout => \GRLFPC20.R.I.EXEC_0_0_G1_0_I_0_0\,
dataa => \GRLFPC20.R.I.EXEC\,
datab => \GRLFPC20.UN1_FPCI_22_X\,
datac => \GRLFPC20.R.I.RDD_0_0_G1_0_574_I_0\,
datad => \GRLFPC20.V.I.EXEC_0_SQMUXA\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110110110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(5),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(6));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_ENTRYPOINT_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT_0\);
GRLFPC20_UN1_MOV_1_SQMUXA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000010000000")
port map (
combout => \GRLFPC20.UN1_MOV_1_SQMUXA_0\,
dataa => \GRLFPC20.COMB.FPDECODE.RDD4_0_A2_0_X\,
datab => \GRLFPC20.MOV_2_SQMUXA_2\,
datac => \GRLFPC20.COMB.FPDECODE.FPOP2_0_A2\,
datad => \GRLFPC20.COMB.FPDECODE.RDD5_0_A3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_EXPBREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\);
GRLFPC20_R_A_MOV_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC20.R.A.MOV_0_0_G1\,
dataa => N_48,
datab => N_49,
datac => \GRLFPC20.R.A.MOV_0_0_G1_3\,
datad => \GRLFPC20.R.A.MOV_0_0_G1_0_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0\,
dataa => N_51,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_5__G0\,
dataa => N_48,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_5__G0_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIS3A83_370_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010110111010010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_0_A3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(370),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_2\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_2_I_O3\);
\GRLFPC20_R_FSR_FTT_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000000000000")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_1__G2_0_624_I\,
dataa => \GRLFPC20.R.X.FPOP\,
datab => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_A6_1_0\,
datac => \GRLFPC20.R.FSR.FTT_1_0_1__G2_0_624_I_1\,
datad => \GRLFPC20.COMB.UN1_MEXC_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_14\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_15\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.NOTAM2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_27\);
\GRLFPC20_R_FSR_FTT_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010001100")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I\,
dataa => \GRLFPC20.R.I.EXC\(5),
datab => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_1\,
datac => \GRLFPC20.COMB.UN1_MEXC_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_7__G0\,
dataa => N_55,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOINSTANDNOEXC_41_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_7__G0_0\);
GRLFPC20_WREN2_1_SQMUXA_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC20.WREN2_1_SQMUXA_1\,
dataa => N_351,
datab => N_352,
datac => \GRLFPC20.WREN1_0_SQMUXA_1_X\,
datad => \GRLFPC20.WREN2_1_SQMUXA_1_1_X\);
GRLFPC20_WREN2_2_SQMUXA_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.WREN2_2_SQMUXA_1\,
dataa => N_339,
datab => \GRLFPC20.R.X.AFSR\,
datac => \GRLFPC20.R.X.LD\,
datad => \GRLFPC20.WREN2_1_SQMUXA_1_1_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001100000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(12),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(13),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(14),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(56),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(27),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(40),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(42),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(44),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(48),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(50),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(51),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(49),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(11),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(21),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(23),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(24),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(25),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(26),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(28),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(29),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(37),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(38),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(39),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(41),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(17),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(18),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(20),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(19),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_A_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(21),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_A_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(47),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(51),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_A_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(45),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_375_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_375__G0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_375__G0_A\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_375_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_375__G0_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_A_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16_A\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(54),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(15),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(14));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1_RNISEO81: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_SUM2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(53),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_113_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(113),
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(113),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_A\(113));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_A_113_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011101000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_A\(113),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(113));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110001010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
GRLFPC20_RS1V_0_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.RS1V_0_SQMUXA\,
dataa => N_74,
datab => N_73,
datac => \GRLFPC20.RS1V_0_SQMUXA_A\,
datad => \GRLFPC20.RS1D_CNST_0_A2_2_X\);
GRLFPC20_RS1V_0_SQMUXA_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000001")
port map (
combout => \GRLFPC20.RS1V_0_SQMUXA_A\,
dataa => N_65,
datab => N_66,
datac => N_62,
datad => N_63);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI3UAN2_370_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001011010010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SUM_I\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(370),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_2_I_O3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN4_STKOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN4_STKOUT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN6_NOTPROP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN2_MIXOIN_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111100001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(371),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_A\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN2_MIXOIN_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011100010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_A\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(43),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110001010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_0_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110001010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_1_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_WQSTSETS_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_WQSTSETS\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN11_WQSTSETS_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(46),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(45));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1_RNICMUB1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN14_CONDITIONAL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN14_CONDITIONAL\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_OPREXCSHFT_UN3_OPREXC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.OPREXCSHFT.UN3_OPREXC\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_4\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_5\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTBZERODENORM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN2_DIVMULTV_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(0));
GRLFPC20_R_I_EXEC_RNO_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010001100")
port map (
combout => \GRLFPC20.R.I.EXEC_0_0_G1_0_I_A8_0\,
dataa => \GRLFPC20.R.I.EXC\(5),
datab => \GRLFPC20.R.I.V\,
datac => \GRLFPC20.COMB.UN1_MEXC_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_16\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(29),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_7__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000010110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_5__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSAMPLEDWAIT\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIIEAL1_315_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110100001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(373),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(315),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN1_NOTPROP_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_NE_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011111111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_NE_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_11_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_12\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_NOTSTICKYINFORSR_2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000100110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.NOTSTICKYINFORSR_2_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN40_SHDVAR\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_RNIRJCN1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM1_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_1_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(1));
\GRLFPC20_R_FSR_FTT_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100000")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_1\,
dataa => \GRLFPC20.R.I.EXEC\,
datab => \GRLFPC20.R.X.FPOP\,
datac => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_0_X\,
datad => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_A6_1_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_16\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_17\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_23\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_24\);
GRLFPC20_COMB_RSDECODE_RS1V2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.COMB.RSDECODE.RS1V2_0\,
dataa => N_52,
datab => N_49,
datac => \GRLFPC20.COMB.RSDECODE.RS1V2_0_A\,
datad => \GRLFPC20.COMB.RSDECODE.UN1_FPCI_0_X\);
GRLFPC20_COMB_RSDECODE_RS1V2_0_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111100000000")
port map (
combout => \GRLFPC20.COMB.RSDECODE.RS1V2_0_A\,
dataa => N_51,
datab => N_50,
datac => N_53,
datad => N_48);
GRLFPC20_COMB_RDD_1_M14_0_A2_0_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100000000000")
port map (
combout => \GRLFPC20.COMB.RDD_1.M14_0_A2_0_0\,
dataa => N_54,
datab => N_55,
datac => N_49,
datad => \GRLFPC20.COMB.RDD_1.M14_0_A2_0_0_A\);
GRLFPC20_COMB_RDD_1_M14_0_A2_0_0_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100100010")
port map (
combout => \GRLFPC20.COMB.RDD_1.M14_0_A2_0_0_A\,
dataa => N_51,
datab => N_50,
datac => N_48,
datad => N_49);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_115_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(115),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(115),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(115),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(115));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI2TFQ_368_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010110111010010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_SUM0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_V\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_EXTEND_TEMP_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1\(1));
GRLFPC20_WREN1_1_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC20.WREN1_1_SQMUXA\,
dataa => \GRLFPC20.WREN1_1_SQMUXA_1\,
datab => \GRLFPC20.WREN1_0_SQMUXA_1_X\,
datac => \GRLFPC20.COMB.UN1_R.I.EXC\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001011010010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI16741_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010101101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_57_SUM0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN26_NOTBINFNAN_4_RNID14F1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_4\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTBINFNAN\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_0\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIA2JO1_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_A\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIGPIQ_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001001110010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_A\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNI1GSQ1_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20_A\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNI7RGD1_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000111110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.TEMP_20_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(71),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(74),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(72));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN4_NOTAINFNAN_RNIQ7TU1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111011100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_4\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTAINFNAN\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_0\(3));
GRLFPC20_ANNULFPU_0_SQMUXA_X_RNIPKTE1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101111")
port map (
combout => \GRLFPC20.ANNULRES_1_SQMUXA\,
dataa => \GRLFPC20.R.X.FPOP\,
datab => \GRLFPC20.R.I.EXEC\,
datac => \GRLFPC20.ANNULFPU_0_SQMUXA_X\,
datad => \GRLFPC20.ANNULRES_1_SQMUXA_A\);
GRLFPC20_ANNULFPU_0_SQMUXA_1_X_RNIBSDG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001100010000")
port map (
combout => \GRLFPC20.ANNULRES_1_SQMUXA_A\,
dataa => \GRLFPC20.R.E.FPOP\,
datab => \GRLFPC20.R.M.FPOP\,
datac => \GRLFPC20.ANNULFPU_0_SQMUXA_2_X\,
datad => \GRLFPC20.ANNULFPU_0_SQMUXA_1_X\);
GRLFPC20_R_A_ST_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.R.A.ST_0_0_G1\,
dataa => \GRLFPC20.N_1243_I_0_A2_1_X\,
datab => \GRLFPC20.COMB.FPDECODE.ST_0_A2\,
datac => CPO_EXCZ,
datad => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I_948_X\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_UN1_ENTRYPOINT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_ENTRYPOINT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_RNIRCSB2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_RNIRCSB2_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_RNIRCSB2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_RNIRCSB2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_RNIRCSB2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN25_NOTXZYFROMD_RNIM5803: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_1_A\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNITOR11_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_1_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN25_NOTXZYFROMD_RNIP8803: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011000110100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_0_A\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIVQR11_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5_0_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN3_NOTXZYFROMD_RNIQ9CH3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000001110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_1_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_CI_114_1_SUM_5_0_A2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010101101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_114_1.SUM_5_0_A2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_RNI9HRN_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010101101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_SUM0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN7_SHDVAR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN7_SHDVAR\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(57));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_38: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_38\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(38));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_37: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_37\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(37));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_35: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_35\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_42: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000111100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_142_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(142),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(142),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(142));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1_RNIIRGN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_AXB0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_172_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_172__G0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLCREGXZ.UN1_INFORCREGDB\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_172__G0_0_M3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.QUOBITS\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_T_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001110110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_T_3\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(377),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.NOTDIVC\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.NOTDIVC\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_R_I_EXC_RNO_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000011100010")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_3__G0\,
dataa => \GRLFPC20.R.I.EXC\(3),
datab => \GRLFPC20.COMB.UN2_HOLDN\,
datac => \GRLFPC20.R.I.EXC_2_0_3__G3\,
datad => \GRLFPC20.COMB.UN19_IUEXEC\);
GRLFPC20_COMB_FPDECODE_RDD3_TZ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.COMB.FPDECODE.RDD3_TZ\,
dataa => N_49,
datab => N_48,
datac => N_51,
datad => \GRLFPC20.COMB.FPDECODE.RDD3_TZ_A\);
GRLFPC20_COMB_FPDECODE_RDD3_TZ_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001111101111")
port map (
combout => \GRLFPC20.COMB.FPDECODE.RDD3_TZ_A\,
dataa => N_53,
datab => N_50,
datac => \GRLFPC20.COMB.FPDECODE.UN1_FPCI_7_1_X\,
datad => \GRLFPC20.COMB.FPDECODE.UN1_FPCI_0_7_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(43));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_43: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_RNIDCD52_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_0\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_RNIDCD52_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN10_NOTPROP_0_2_I_O3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_0\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_UN53_SCTRL_NEW: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.UN53_SCTRL_NEW\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_NORMDETECT_NOTSLFROMNORM_17_3_0__M3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110100011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN30_CONDITIONAL_M5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111100010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M2_E_4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M2_E_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M5_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN30_CONDITIONAL_M5_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010101010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M5_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_NORMDETECT_NOTSLFROMNORM_17_3_0__M2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110100011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_NORMDETECT_NOTSLFROMNORM_17_3_0__M4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001110100011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.NORMDETECT.NOTSLFROMNORM_17_3_0_.M4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_235_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(235),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(235),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(235),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_EXPAREGLOADEN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100111011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_234_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(234),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(234),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(234),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_236_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(236),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(236),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(236),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.RESULT\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\);
GRLFPC20_COMB_V_I_EXEC_5_IV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC20.COMB.V.I.EXEC_5_IV\,
dataa => \GRLFPC20.R.I.EXEC\,
datab => \GRLFPC20.UN1_FPCI_22_X\,
datac => \GRLFPC20.V.I.EXEC_0_SQMUXA\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_10\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN36_STKGEN_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111101110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN36_STKGEN_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN11_WQSTSETS_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110001010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN11_WQSTSETS_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN4_NOTSHIFTCOUNT1_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TEMP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_ENTRYPOINT_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.ENTRYPOINT_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.ENTRYSHFT.S_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_EXTEND_TEMP_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1_A\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_EXTEND_TEMP_1_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001101011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1_A\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(230),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_RNO_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_1_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(218),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_RNO_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(220),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_RNO_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3_E_0_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(219),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN3_NOTBZERODENORM_RNI8BNJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010100010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_0\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTBZERODENORM\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN3_NOTAZERODENORM_0_RNIO7OP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_0\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM_0\);
GRLFPC20_WREN1_1_SQMUXA_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.WREN1_1_SQMUXA_1\,
dataa => N_351,
datab => N_352,
datac => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datad => \GRLFPC20.R.X.SEQERR\(0));
GRLFPC20_COMB_RDD_1_M14_0_A2_0_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001000000000")
port map (
combout => \GRLFPC20.COMB.RDD_1.M14_0_A2_0_1\,
dataa => N_49,
datab => N_48,
datac => N_54,
datad => \GRLFPC20.COMB.FPDECODE.RDD4_0_A2_0_X\);
GRLFPC20_COMB_FPDECODE_FPOP8_I_O3_X_RNI8EF33: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.R.A.AFQ_0_0_G1_0\,
dataa => N_65,
datab => N_66,
datac => N_63,
datad => \GRLFPC20.R.A.AFQ_0_0_G1_0_3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M14S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14S2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8S2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11S4\);
GRLFPC20_COMB_RSDECODE_UN1_FPCI_0_X_RNIGOBD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.R.A.RS1D_0_0_G4\,
dataa => N_51,
datab => N_53,
datac => \GRLFPC20.R.A.RS1D_0_0_G4_1_X\,
datad => \GRLFPC20.COMB.RSDECODE.UN1_FPCI_0_X\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_DPATH_NEW_7_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA_0\,
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\);
GRLFPC20_RS2_0_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.RS2_0_SQMUXA\,
dataa => N_65,
datab => N_63,
datac => \GRLFPC20.RS2_0_SQMUXA_0_X\,
datad => \GRLFPC20.COMB.V.A.RF1REN_1_0_650_A2_3_X\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_COUNTSUCCESSIVEZERO18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_10\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(12));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000011101111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(10));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN3_NOTAZERODENORM_0_RNIVK541: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_4\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_5\(5),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM_0\);
GRLFPC20_COMB_UN9_CCV_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000111")
port map (
combout => CPO_CCVZ,
dataa => N_269,
datab => \GRLFPC20.R.M.FPOP\,
datac => \GRLFPC20.COMB.UN9_CCV_0_0\,
datad => \GRLFPC20.COMB.UN9_CCV_0_1\);
GRLFPC20_COMB_UN19_IUEXEC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.COMB.UN19_IUEXEC\,
dataa => \GRLFPC20.R.MK.BUSY2\,
datab => \GRLFPC20.R.MK.BUSY\,
datac => \GRLFPC20.FPI.LDOP_2\,
datad => \GRLFPC20.COMB.LOCKGEN.DEPCHECK\);
\GRLFPC20_R_I_EXC_RNO_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010101000")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_4__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STATUS\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DECODESTATUS.UN7_STATUS\,
datad => \GRLFPC20.COMB.UN2_HOLDN\);
GRLFPC20_COMB_UN1_MEXC_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000000000000")
port map (
combout => \GRLFPC20.COMB.UN1_MEXC_1\,
dataa => \GRLFPC20.R.FSR.TEM\(1),
datab => \GRLFPC20.R.I.EXC\(1),
datac => \GRLFPC20.COMB.UN1_MEXC_1_0\,
datad => \GRLFPC20.COMB.UN1_MEXC_1_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_UN10_S_MOV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_UN1_ENTRYPOINT_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110100111111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_UN1_ENTRYPOINT_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001101100101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN1_S_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_EXTEND_TEMP_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111110101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI8QPI_228_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(228),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI7PPI_227_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(227),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI6OPI_226_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(226),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI5NPI_225_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(225),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI4MPI_224_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(224),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI3LPI_223_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(223),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI2KPI_222_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(222),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_4\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(7),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M4_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIV1H32_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101111111110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0_A2_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_32_0_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTNULLEXC\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77));
GRLFPC20_R_I_RDD_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000010100000")
port map (
combout => \GRLFPC20.R.I.RDD_0_0_G1_0_574_I\,
dataa => \GRLFPC20.R.I.RDD\,
datab => \GRLFPC20.R.X.RDD\(0),
datac => \GRLFPC20.R.I.RDD_0_0_G1_0_574_I_0\,
datad => \GRLFPC20.V.I.EXEC_0_SQMUXA\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_SIGNRESULT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.SIGNRESULT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(23),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.UN1_GRFPUS\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2_RNI1EP4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_2_RNI0NR1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_1_RNIUVTE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_3_RNIV80C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_2_RNITH29: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1_RNI49P2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_RNIJIT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1_RNI2RTC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3_RNI340A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3_RNI2D27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3_RNI1M44: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2_RNIVU61: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_RNIDKDD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_1_RNISGBB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_1_RNIRPD8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_RNIJH8E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3_RNI4Q6F: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_1_RNI139C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2_RNI0LD6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_2_RNIVTF3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_3_RNIV6I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2_RNITFKD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2_RNISOMA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3_RNIS1P7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_2_RNI3PF1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_1_RNI12IE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1_RNI0BKB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_RNIDI38: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2_RNITETF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3_RNITNVC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_RNIH5P7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_RNIGG6F: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_3_RNI1JVA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2_RNIVR18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_RNIDHE5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2_RNITD62: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3_RNIR8D9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3_RNIQHF6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2_RNIH597: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2_RNIGEB4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3_RNIGND1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_RNITCJ9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3_RNIE9IB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3_RNIDIK8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_RNIQDRF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3_RNIB4P2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_CIN_10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_CIN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.CIN_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_RNIU1IA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_RNITCVH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_RNISNC9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3_RNIM0M4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_RNIKIQE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2_RNIIRSB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1_RNIG4V8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2_RNIGD16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3_RNIGM33: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3_RNIFV5G: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_RNIE88D: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_RNIDHAA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_RNIK814: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1_RNIIH3H: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2_RNIIQ5E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_RNIELC5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_RNIDUE2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_RNIDGJC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2_RNIBPL9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_RNI2JT4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_RNIJPEG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_RNI09O3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2_RNIETN4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1_RNIC6QH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_RNIRVQ8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3_RNICOUB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_RNIPLL7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1_RNIHON2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1_RNIG1QF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_RNIVIG8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_RNIGJU9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2_RNIES07: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_RNIOVDC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_RNIG385: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1_RNIV586: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_RNIEP24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1_RNITNCG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2_RNIT0FD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_RNIBQAA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3_RNIHMJL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_RNI7C1M: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_1_RNIK8HM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_RNI3OMJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_RNI234R: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_2_RNIHCQQ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_RNIGLSN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_2_RNIFUUK: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1_RNIMLLE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2_RNIMUNR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_RNI4CKP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_1_RNIJGSL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_RNI22FO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_RNI1DSF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_RNI0O9N: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_RNIV2NE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1_RNIET7N: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_1_RNID6AK: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_RNIHJES: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_RNIE5JM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_3_RNIM5CD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3_RNILEEQ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_RNIJNGN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_RNI1BIQ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3_RNII9LH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3_RNIHINE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2_RNIFRPR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_2_RNIDDUL: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_RNIBM0J: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1_RNI3AQJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_RNIIR9N: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1_RNI1SUD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3_RNI251R: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_RNIVD3O: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1_RNIUM5L: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_RNITV7I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_RNIT8AF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1_RNIRHCS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_RNIVM43: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.CIN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_UN35_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2_RNI1CB9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_RNI1EHI: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3_RNINT0E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_RNI4BVM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1_RNIH1AI: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_1_RNIGACF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_UN5_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111101110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_UN5_ZERO_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_14_142_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_14\(142),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(144),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.QUOBITS\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3_RNIESA6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_RNIC5DJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1_RNIAEFG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_RNI9NHD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2_RNIIE87: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_1_RNIGNAK: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2_RNIG0DH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_RNIUD7K: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_2_RNIEIHB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_RNICRJ8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1_RNIB4M5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1_RNIADOI: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_RNIP4A9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_RNIOFNG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_RNIIMJ6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_RNIV15A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_3_RNIG8OG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_RNITNV8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_3_RNIEQSA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_3_RNID3V7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_2_RNIBC15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_RNI9L3I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_RNIOE2E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_RNINPF5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1_RNIFUU5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_2_RNIF71J: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3_RNIFG3G: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_2_RNIDP5D: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_3_RNID28A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_RNICBA7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_1_RNI6FJB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2_RNIF6A5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_2_RNIEFCI: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1_RNICOEF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_RNI6ESD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2_RNI6NUA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3_RNIVAOB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_3_RNIUJQ8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_2_RNISSS5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_RNIR5VI: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_RNI9TF5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2_RNIPN3D: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_RNIP06A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1_RNIM987: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_RNI595J: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.2.CI_56_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_UN20_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_RNIP20K: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1_RNI8TEH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_1_RNI76HE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_1_RNIB1HC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1_RNIAAJ9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1_RNI9JL6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(185),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(192),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(202),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(205),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(206),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(208),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(213),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(214),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6_A\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_A_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6_A\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(44),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(175),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(177),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(178),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(181),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(182),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(183),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(184),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(186),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(187),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(189),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(191),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(193),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(194),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(196),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(197),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(198),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(199),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(201),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(203),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(207),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(209),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(210),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(212),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(215),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(216),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101111101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(57),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_A_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_A_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(35),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_46__G2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_21__G2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(41),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_20__G2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_20__G2_A\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_41\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_15\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010100101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_20__G2_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD10_RNIED4Q: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRTOSTICKY\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TEMP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD11\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN12_SRTOSTICKY_3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(190),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(180),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(179),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(176),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(57));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN40_SHDVAR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN40_SHDVAR\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2_0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1_RNIDJ89: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2_RNIFA6C: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_7356\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_3_RNILIAH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.CIN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1_RNIIRCE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.N_1299_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_RNI11A4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.CIN_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3_RNIQ4OH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_RNI9G59: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_RNIRIJ7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_MOV_7_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.MOV_7_SQMUXA\,
dataa => N_62,
datab => N_64,
datac => \GRLFPC20.COMB.FPDECODE.FPOP3_0\,
datad => \GRLFPC20.COMB.V.A.RF1REN_1_0_650_A2_3_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(188),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_RNI52SK: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2_RNINMCS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3_RNIE7HF: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3_RNIL9OH: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_173_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_173__G0_I\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(173),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(56),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(55));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_CIN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2_RNIODQE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_3_RNIASNJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_RNINN5G: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN20_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_UN50_ZERO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2_RNIE4SO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2_RNIFSGP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_RNIPK05: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_RNIAN7E: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1_RNIBE5H: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_RNISJOE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3_RNISVAC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_RNIB794: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_SCTRL_NEW_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_A\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_SCTRL_NEW_A_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_A\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(2),
datab => \GRLFPC20.R.FSR.RD\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(54));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN2_NOTABORTWB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110111001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTNULLEXC\,
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M14_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14S2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M14_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14S2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M14_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14S2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M14_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M14S2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2_1\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(7),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(9),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_EXPYBUS_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_EXPYBUS_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_EXPYBUS_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(240),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(240),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(240),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(241),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(241),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(241),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(242),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(242),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(242),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(238),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(238),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(238),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(244),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(244),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(243),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(243),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(243),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(239),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(239),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(239),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(237),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(237),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(237),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(195),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1_RNIFCA8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3_RNII38B: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100001001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_6_0_67__G3\,
dataa => N_54,
datab => N_62,
datac => N_56,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_1_X\);
GRLFPC20_COMB_LOCKGEN_LOCKI_I_0_0_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100001111")
port map (
combout => \GRLFPC20.COMB.LOCKGEN.LOCKI_I_0_0_A2_0\,
dataa => N_73,
datab => N_74,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.COMB.FPDECODE.ST3_1\);
GRLFPC20_V_FSR_FTT_1_SQMUXA_0_RNIDF1F1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101011111010")
port map (
combout => \GRLFPC20.UN1_FPCI_13\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.AFQ\,
datac => \GRLFPC20.V.FSR.FTT_1_SQMUXA_0\,
datad => \GRLFPC20.COMB.QNE2\);
GRLFPC20_R_X_AFQ_RNI5DJ81: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101110101111")
port map (
combout => \GRLFPC20.UN1_FPCI_2\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.AFQ\,
datac => \GRLFPC20.R.X.SEQERR\(0),
datad => \GRLFPC20.COMB.QNE2\);
GRLFPC20_COMB_RDD_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011110000")
port map (
combout => \GRLFPC20.COMB.RDD_2\,
dataa => \GRLFPC20.COMB.UN1_FPCI_0_X\,
datab => \GRLFPC20.R.X.RDD\(0),
datac => \GRLFPC20.R.I.RDD\,
datad => \GRLFPC20.COMB.UN1_R.I.V_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_6\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(47));
\GRLFPC20_COMB_V_FSR_CEXC_1_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(4),
dataa => \GRLFPC20.R.I.EXC\(4),
datab => \GRLFPC20.R.FSR.TEM\(4),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(4),
datad => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC20_COMB_V_FSR_CEXC_1_2_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(3),
dataa => \GRLFPC20.R.I.EXC\(3),
datab => \GRLFPC20.R.FSR.TEM\(3),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(3),
datad => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC20_COMB_V_FSR_CEXC_1_2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(2),
dataa => \GRLFPC20.R.I.EXC\(2),
datab => \GRLFPC20.R.FSR.TEM\(2),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(2),
datad => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC20_COMB_V_FSR_CEXC_1_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(1),
dataa => \GRLFPC20.R.I.EXC\(1),
datab => \GRLFPC20.R.FSR.TEM\(1),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(1),
datad => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M2\);
\GRLFPC20_COMB_V_FSR_CEXC_1_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001111")
port map (
combout => \GRLFPC20.COMB.V.FSR.CEXC_1_2\(0),
dataa => \GRLFPC20.R.I.EXC\(0),
datab => \GRLFPC20.R.FSR.TEM\(0),
datac => \GRLFPC20.COMB.V.FSR.CEXC_1_2_A_X\(0),
datad => \GRLFPC20.COMB.V.FSR.CEXC_1_SN_M2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_RNIEELJ: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_2_RNIQ947: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_RNIAJBE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3_RNISQEP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010110011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0_A\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(30),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(211),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(204),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_NOTSRRES_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_NOTSRRES_0\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3_RNIKO7L: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_2_RNIKF5O: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_2_RNIHDHO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3_RNIJ4FR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN35_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_RNIUUI2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_RNIVJ5B: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN50_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_2_RNIVSO5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1_RNIVJM8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.UN5_ZERO\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_SCTRL_39_IV_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL_I_M_1\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.UN4_TEMP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_EXTEND_TEMP_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.EXTEND.TEMP_1\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN26_XZYBUSLSBS\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_UN3_S_SQRT_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_24\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_23: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_23\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_18\);
\GRLFPC20_R_FSR_FTT_RNO_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000000000")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_1__G2_0_624_I_1\,
dataa => \GRLFPC20.R.I.EXEC\,
datab => \GRLFPC20.R.X.FPOP\,
datac => \GRLFPC20.R.I.EXC\(5),
datad => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_0_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIJFAQ_229_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M4_1_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(229),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_UN23_EXPXBUS_11_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.UN23_EXPXBUS_11_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(11));
\GRLFPC20_R_X_SEQERR_RNI435M_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I_A6_1_0\,
dataa => N_354,
datab => N_353,
datac => N_4,
datad => \GRLFPC20.R.X.SEQERR\(0));
GRLFPC20_R_A_MOV_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.R.A.MOV_0_0_G1_3\,
dataa => N_55,
datab => N_56,
datac => \GRLFPC20.R.A.MOV_0_0_G1_1_X\,
datad => \GRLFPC20.COMB.FPDECODE.RDD5_3_0_A2_X\);
GRLFPC20_MOV_2_SQMUXA_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC20.MOV_2_SQMUXA_2\,
dataa => N_55,
datab => N_56,
datac => N_52,
datad => \GRLFPC20.COMB.FPDECODE.RDD4_0_A2_X\);
GRLFPC20_COMB_FPDECODE_FPOP8_I_O3_X_RNI13GO1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC20.R.A.AFQ_0_0_G1_0_3\,
dataa => N_64,
datab => N_62,
datac => N_67,
datad => \GRLFPC20.COMB.FPDECODE.FPOP8_I_O3_X\);
GRLFPC20_COMB_FPDECODE_RDD5_0_A3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.RDD5_0_A3\,
dataa => N_49,
datab => N_48,
datac => \GRLFPC20.COMB.FPDECODE.RDD5_3_0_A2_X\,
datad => \GRLFPC20.COMB.RSDECODE.UN1_FPCI_0_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_52_RNIJOM31\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_9__G4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_52\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN17_SHDVAR: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_A\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN17_SHDVAR_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN3_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD_A\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN3_NOTXZYFROMD_A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD_A\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111100011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN33_PCTRL_NEW_I_0_G0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(61),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M13_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11S4\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLAREGXZ_UN5_XZAREGLOADEN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLAREGXZ.UN5_XZAREGLOADEN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datad => \GRLFPC20.FPI.LDOP\);
GRLFPC20_COMB_LOCKGEN_DEPCHECK: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111111")
port map (
combout => \GRLFPC20.COMB.LOCKGEN.DEPCHECK\,
dataa => \GRLFPC20.R.M.FPOP\,
datab => \GRLFPC20.R.X.FPOP\,
datac => \GRLFPC20.R.A.FPOP\,
datad => \GRLFPC20.ANNULRES_0_SQMUXA_12_1\);
GRLFPC20_COMB_UN2_HOLDN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC20.COMB.UN2_HOLDN\,
dataa => \GRLFPC20.COMB.UN3_HOLDN_X\,
datab => N_3,
datac => \GRLFPC20.R.A.FPOP\,
datad => \GRLFPC20.R.A.MOV\);
\GRLFPC20_R_I_EXC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC20.R.I.EXC_0\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DECODESTATUS.UN7_STATUS\,
datad => \GRLFPC20.COMB.UN2_HOLDN\);
\GRLFPC20_R_I_EXC_RNO_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_3__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
datad => \GRLFPC20.COMB.UN2_HOLDN\);
GRLFPC20_COMB_FPDECODE_FPOP2_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.FPOP2_0_A2\,
dataa => N_64,
datab => N_66,
datac => \GRLFPC20.COMB.RDD_1.M10_2_0_A2_X\,
datad => \GRLFPC20.COMB.FPDECODE.FPOP2_0_O2_X\);
GRLFPC20_COMB_LOCK_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => CPO_LDLOCKZ,
dataa => N_77,
datab => \GRLFPC20.R.STATE\(0),
datac => \GRLFPC20.R.STATE\(1),
datad => \GRLFPC20.COMB.LOCK_1_1_X\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_S_CMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN3_NOTXZYFROMD_RNIUMVM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN3_NOTXZYFROMD_RNIV28P: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN3_NOTXZYFROMD_RNI477P: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_3_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIK3451_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011111111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD12_RNI5OTA1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_E\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD12\,
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
GRLFPC20_R_A_MOV_RNIOME21: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000101010101010")
port map (
combout => \GRLFPC20.R.I.RDD_0_0_G1_0_574_I_0\,
dataa => N_1,
datab => \GRLFPC20.COMB.UN3_HOLDN_X\,
datac => \GRLFPC20.R.A.FPOP\,
datad => \GRLFPC20.R.A.MOV\);
GRLFPC20_V_FSR_AEXC_1_SQMUXA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111100000000")
port map (
combout => \GRLFPC20.V.FSR.AEXC_1_SQMUXA_0\,
dataa => N_389,
datab => N_388,
datac => N_390,
datad => \GRLFPC20.V.FSR.NONSTD_0_SQMUXA_2_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_0_A2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_0_A2\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_41__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_A\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_A_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_A\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_45\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_RNIRQQ9_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_TEMP_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_RNIP5VG_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.TEMP_2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110110001101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_0\(4));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_57: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(57));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN18_XZXBUS_31: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN18_XZXBUS_31\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(31));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN4_NOTBINFNAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTBINFNAN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_115_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(115),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.ROMXZSL2FROMC\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(61),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(61));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(62));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(63),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(63));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(64),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(64));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(65),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(65));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(66),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(66));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(67),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(67));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(68),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(68));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(69),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(69));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(70),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(70));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(71),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(71));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(72),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(72));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(73),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(73));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(74),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(74));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(76),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(76));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(77),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(77));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(78),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(78));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(79),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(79));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(80),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(80));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(81),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(81));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(82),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(82));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(126),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(128),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(129),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(132),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(16));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_GRFPUF_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELINITREMBIT_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_0_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_A\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_0_A_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_A\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_A\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_0_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_0_A\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(120),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(122),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(6));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_142_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(142),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_A_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3_A\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(121),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(124),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(127),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(130),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(133),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(135),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(136),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(138),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(140),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1_X\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1_X\(25));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(125),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(134),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(137),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(139),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1_X\(23));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.8.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.37.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.19.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.38.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.23.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.6.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.9.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.39.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.24.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.18.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.34.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.40.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.41.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.42.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.10.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.29.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.30.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.31.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.16.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.7.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.49.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.44.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.28.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.45.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.46.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.5.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.43.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.33.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.15.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.17.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.4.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.50.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(62),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(62));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_0_A2\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_61\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.ENTRYSHFT.S_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(62));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(61),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_58\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.ENTRYSHFT.S_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(61));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010111000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(60),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_59\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_I_O2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(60));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(59),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_I_O2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010111000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_49\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_I_O2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.ENTRYSHFT.S_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_A\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_A_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_A\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(39),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_A\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_A_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111000111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_A\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_16\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN6_S_0_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN6_S_0_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_20\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_19\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN6_S_0_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_0_A2\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(12),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M5S4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_41__G4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_9__G3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_112__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(112));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_109__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(109));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_107__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(107));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_106__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(106));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_105__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(105));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_104__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(104));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_103__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(103));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_100__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(100));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_99__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(99));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_98__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(98));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_97__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(97));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_96__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(96));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_94__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(94));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_92__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(92));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_90__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(90));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_89__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(89));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_88__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(88));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_86__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(86));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_84__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_141_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(141),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN23_XZROUNDOUT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN23_XZROUNDOUT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(131),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.53.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_54_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.54.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(53));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_55_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.55.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_111__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(111));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_172_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_172__G0_0_M3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_171_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(171),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_23_113_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110001001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(113),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_95__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(95));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_108__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(108));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_110__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(110));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.3.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.1.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.2.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.32.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.48.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.47.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(123),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIDLA61_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000011100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110101011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(49));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIK8201_372_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN1_NOTPROP_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(372),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(114),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.ROMXZSL2FROMC\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_91__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(91));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULLSBLOGIC_STCKYPAIR_UN4_STKOUT_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101001011010010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULLSBLOGIC.STCKYPAIR.UN6_NOTPROP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(371),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_101__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(101));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_102__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(102));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.22.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.11.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.14.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.12.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.13.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_SCTRL_NEW_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011101000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLAREGEXP_EXPAREGLOADEN_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLAREGEXP.EXPAREGLOADEN_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD12\,
datac => \GRLFPC20.FPI.LDOP\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_6_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101101000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_6\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UPDATE_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(71),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(72),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M12_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M12_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M13_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11S4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M13_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11S4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M13_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M13\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8S2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11S4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M12_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000111110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M12\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100011111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_26_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_26\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2_1\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_EXPYBUS_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_EXPYBUS_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(240),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(240),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(241),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(241),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(242),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(242),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_235_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(235),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP2_X\(61),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(238),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(238),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(244),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_233_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(233),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_A\(233),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_A_233_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100111101111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_A\(233),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD11\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M11S4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11S4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_236_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(236),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP2_X\(60),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_234_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(234),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datac => \GRLFPC20.FPI.OP2_X\(62),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(243),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(243),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(239),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(239),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(237),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(237),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_232_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110000001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(232),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(232),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(232));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN4_NOTAINFNAN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN4_NOTAINFNAN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.36.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.35.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_GRFPUF_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELINITREMBIT_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_GRFPUF_0_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELINITREMBIT_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_GRFPUF_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000011011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELINITREMBIT_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELINITREMBIT_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIVA8D1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_37\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51));
GRLFPC20_COMB_UN1_FPCI_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001000100010")
port map (
combout => \GRLFPC20.COMB.UN1_FPCI_4\,
dataa => \GRLFPC20.R.A.RS2\(0),
datab => \GRLFPC20.R.A.RS2D\,
datac => \GRLFPC20.R.A.RS1D\,
datad => \GRLFPC20.COMB.UN1_FPCI_0_1_X\);
GRLFPC20_COMB_UN1_R_A_RS1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110000")
port map (
combout => \GRLFPC20.COMB.UN1_R.A.RS1_1\,
dataa => N_145,
datab => \GRLFPC20.R.A.ST\,
datac => \GRLFPC20.R.A.RS1\(0),
datad => \GRLFPC20.R.A.RS1D\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN3_INEXACT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000001110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN3_INEXACT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.NOTAM2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_0__G0_0\,
dataa => N_50,
datab => N_54,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_0__G0_0_A3_0_X\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MAPMULXFF.UN4_UNIMPMAP_1_X\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_5_0_1__G0\,
dataa => N_55,
datab => N_52,
datac => N_54,
datad => N_50);
GRLFPC20_COMB_RDD_1_M14_0_A2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.COMB.RDD_1.M14_0_A2_1\,
dataa => N_66,
datab => N_64,
datac => \GRLFPC20.COMB.FPDECODE.FPOP2_0_O2_X\,
datad => \GRLFPC20.COMB.FPDECODE.FPOP8_I_O3_X\);
GRLFPC20_COMB_V_A_AFSR_1_5_0_O2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC20.COMB.V.A.AFSR_1_5_0_O2_1\,
dataa => N_62,
datab => N_63,
datac => N_64,
datad => \GRLFPC20.COMB.FPDECODE.FPOP2_0_O2_X\);
GRLFPC20_COMB_FPDECODE_ST_0_A2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.ST_0_A2\,
dataa => N_65,
datab => N_66,
datac => \GRLFPC20.RS1D_CNST_0_A2_2_X\,
datad => \GRLFPC20.COMB.FPDECODE.FPOP8_I_O3_X\);
GRLFPC20_V_I_EXEC_0_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC20.V.I.EXEC_0_SQMUXA\,
dataa => N_354,
datab => N_353,
datac => N_4,
datad => \GRLFPC20.R.X.FPOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_7_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_14_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN8_TEMP_U_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111100000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_U\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_2\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN15_XZROUNDOUT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_85__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_93__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(93));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.20.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.21.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_A_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_A\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M3_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(83),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(83));
GRLFPC20_WRADDR_1_SQMUXA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101010101")
port map (
combout => \GRLFPC20.WRADDR_1_SQMUXA\,
dataa => \GRLFPC20.WRADDR_0_SQMUXA_0_X\,
datab => \GRLFPC20.R.I.EXEC\,
datac => \GRLFPC20.R.I.V\,
datad => \GRLFPC20.R.X.FPOP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100011011000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNO_0_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_87__G1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(87));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.52.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.25.TRFWWBASICCELL.TEMP2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.51.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.26.TRFWWBASICCELL.TEMP2_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101101000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.27.TRFWWBASICCELL.TEMP2_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(119),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIHQJ91_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
datac => \GRLFPC20.FPI.LDOP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_CHECKOVANDDENORM_UN13_NOTPOSSIBLEOV_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.CHECKOVANDDENORM.UN13_NOTPOSSIBLEOV_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIHQJ91_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_0_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
datac => \GRLFPC20.FPI.LDOP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN30_CONDITIONAL_M2_E_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M2_E_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD3\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD6\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN30_CONDITIONAL_M2_E_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN30_CONDITIONAL_M2_E_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNI3F121_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_1\(77),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(46));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN17_SHDVAR_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN17_SHDVAR_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(2));
GRLFPC20_R_A_AFSR_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.R.A.AFSR_0_0_G1_1_0\,
dataa => N_62,
datab => N_67,
datac => N_63,
datad => N_65);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_UN10_S_MOV_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN10_S_MOV_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN12_SRTOSTICKY_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN12_SRTOSTICKY_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD6\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD9\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_18\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_17\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_16\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_15\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_13: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35));
GRLFPC20_COMB_UN1_MEXC_1_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC20.COMB.UN1_MEXC_1_1\,
dataa => \GRLFPC20.R.FSR.TEM\(3),
datab => \GRLFPC20.R.I.EXC\(3),
datac => \GRLFPC20.R.FSR.TEM\(0),
datad => \GRLFPC20.R.I.EXC\(0));
GRLFPC20_COMB_UN1_MEXC_1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101110111")
port map (
combout => \GRLFPC20.COMB.UN1_MEXC_1_0\,
dataa => \GRLFPC20.R.FSR.TEM\(4),
datab => \GRLFPC20.R.I.EXC\(4),
datac => \GRLFPC20.R.FSR.TEM\(2),
datad => \GRLFPC20.R.I.EXC\(2));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_COUNTSUCCESSIVEZERO18_11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_COUNTSUCCESSIVEZERO18_10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_COUNTSUCCESSIVEZERO18_9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_COUNTSUCCESSIVEZERO18_8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_COUNTSUCCESSIVEZERO18_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNINA99_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_5\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIOA89_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_4\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN26_NOTBINFNAN_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN26_NOTBINFNAN_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTBINFNAN_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN26_NOTAINFNAN_5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN26_NOTAINFNAN_4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN26_NOTAINFNAN_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_OPREXCSHFT_UN3_OPREXC_RNO_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_5\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_OPREXCSHFT_UN3_OPREXC_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS_4\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252));
GRLFPC20_V_FSR_FTT_1_SQMUXA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110100001101")
port map (
combout => \GRLFPC20.V.FSR.FTT_1_SQMUXA_0\,
dataa => \GRLFPC20.R.X.AFSR\,
datab => \GRLFPC20.R.X.LD\,
datac => \GRLFPC20.R.X.SEQERR\(0));
GRLFPC20_COMB_UN9_CCV_0_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC20.COMB.UN9_CCV_0_1\,
dataa => N_338,
datab => \GRLFPC20.R.X.FPOP\,
datac => \GRLFPC20.R.I.EXEC\,
datad => \GRLFPC20.R.I.INST\(19));
GRLFPC20_COMB_UN9_CCV_0_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC20.COMB.UN9_CCV_0_0\,
dataa => N_200,
datab => \GRLFPC20.R.E.FPOP\,
datac => \GRLFPC20.R.X.AFSR\,
datad => \GRLFPC20.R.X.LD\);
GRLFPC20_COMB_FPDECODE_RDD3_TZ_A_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.UN1_FPCI_0_7_2\,
dataa => N_54,
datab => N_55,
datac => N_52,
datad => N_53);
GRLFPC20_COMB_FPDECODE_FPOP3_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.FPOP3_0\,
dataa => N_66,
datab => N_67,
datac => N_63,
datad => N_65);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD56_RNI5SGF1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WQSTSETS\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_4_0_2__G0\,
dataa => N_54,
datab => N_50,
datac => N_55,
datad => N_52);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1_520\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(2),
datab => \GRLFPC20.R.FSR.RD\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_WQSCTRL_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.WQSCTRL\(68),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD12\,
datac => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIDLA61_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN3_NOTBZERODENORM: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTBZERODENORM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_4_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111101111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51));
GRLFPC20_COMB_V_A_LD_1_0_A2_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.COMB.V.A.LD_1_0_A2_0\,
dataa => \GRLFPC20.R.M.LD\,
datab => \GRLFPC20.R.X.LD\,
datac => \GRLFPC20.R.A.LD\,
datad => \GRLFPC20.R.E.LD\);
GRLFPC20_FPI_LDOP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111111101")
port map (
combout => \GRLFPC20.FPI.LDOP\,
dataa => N_1,
datab => \GRLFPC20.R.MK.LDOP\,
datac => \GRLFPC20.R.MK.RST\,
datad => \GRLFPC20.R.MK.RST2\);
GRLFPC20_COMB_UN1_R_I_V_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.COMB.UN1_R.I.V_0\,
dataa => \GRLFPC20.R.I.EXEC\,
datab => \GRLFPC20.R.I.V\,
datac => \GRLFPC20.R.X.FPOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNI8Q721_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI5IJD1_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.NOTAM2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_1_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIAR1O_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0_A2_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0_REP2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN15_NOTXZYFROMD_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN15_NOTXZYFROMD_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_RNDMODESELECT_UN17_U_RDN: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.UN17_U_RDN\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
datab => \GRLFPC20.R.FSR.RD\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.UN17_U_RDN_I_0_503_I_A2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
datab => \GRLFPC20.R.FSR.RD\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010001010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_19\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_0_A2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_0_A2\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(310),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(309),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(308),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(307),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(306),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(305),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(304),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(303),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(302),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(300),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(297),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(296),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(294),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(292),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(290),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(289),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(288),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(286),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(284),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(282),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(280),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(279),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(275),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(274),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(272),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(271),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(270),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(269),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(268),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(266),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(264),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(263),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(262),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(261),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(260),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_SHIFT_4_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_4\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_SHIFT_3_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_3\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIVCHI1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(298),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(295),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(291),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(285),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(281),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(276),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_SHIFT_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_1\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_17\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_MULTIPLELOGIC_SHIFT_2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010111001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.MULTIPLELOGIC.SHIFT_2\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(5));
\GRLFPC20_COMB_DBGDATA_4_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(29),
dataa => N_621,
datab => N_685,
datac => N_391,
datad => N_390);
\GRLFPC20_COMB_DBGDATA_4_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111001010")
port map (
combout => CPO_DBG_DATAZ(18),
dataa => N_610,
datab => N_674,
datac => N_391,
datad => N_390);
\GRLFPC20_COMB_DBGDATA_4_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111001010")
port map (
combout => CPO_DBG_DATAZ(17),
dataa => N_609,
datab => N_673,
datac => N_391,
datad => N_390);
\GRLFPC20_COMB_DBGDATA_4_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(21),
dataa => N_613,
datab => N_677,
datac => N_391,
datad => N_390);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(61),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(61));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(62));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(63),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(63));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(64),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(64));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(65),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(65));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(66),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(66));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(67),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(67));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(68),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(68));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(69),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(69));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(70),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(70));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(71),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(71));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(72),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(72));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(73),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(73));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(74),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(74));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(76),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(76));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(77),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(77));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(78),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(78));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(79),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(79));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(80),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(80));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(81),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(81));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(82),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(82));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(84),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(86),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(86));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(88),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(88));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(89),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(89));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(90),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(90));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(92),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(92));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(94),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(94));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(96),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(96));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(97),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(97));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(98),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(98));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(99),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(99));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(100),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(100));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(103),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(103));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(104),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(104));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(105),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(105));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(106),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(106));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(107),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(107));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(109),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(109));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(112),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(112));
\GRLFPC20_COMB_RS1_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110000000")
port map (
combout => \GRLFPC20.COMB.RS1_1\(1),
dataa => N_69,
datab => \GRLFPC20.RS1V_0_SQMUXA\,
datac => \GRLFPC20.COMB.RS1_1_SN_M2_X\,
datad => \GRLFPC20.COMB.RS1_1_0_X\(1));
\GRLFPC20_COMB_V_E_STDATA_1_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(2),
dataa => \GRLFPC20.R.FSR.CEXC\(2),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(34));
\GRLFPC20_COMB_V_E_STDATA_1_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(4),
dataa => \GRLFPC20.R.FSR.CEXC\(4),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(36));
\GRLFPC20_COMB_V_E_STDATA_1_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(5),
dataa => \GRLFPC20.R.FSR.AEXC\(0),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(37));
\GRLFPC20_COMB_V_E_STDATA_1_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(7),
dataa => \GRLFPC20.R.FSR.AEXC\(2),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(39));
\GRLFPC20_COMB_V_E_STDATA_1_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(8),
dataa => \GRLFPC20.R.FSR.AEXC\(3),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(40));
\GRLFPC20_COMB_V_E_STDATA_1_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(10),
dataa => CPO_CCZ(0),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(42));
\GRLFPC20_COMB_V_E_STDATA_1_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(23),
dataa => \GRLFPC20.R.FSR.TEM\(0),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(55));
\GRLFPC20_COMB_V_E_STDATA_1_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(24),
dataa => \GRLFPC20.R.FSR.TEM\(1),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(56));
\GRLFPC20_COMB_V_E_STDATA_1_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(26),
dataa => \GRLFPC20.R.FSR.TEM\(3),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(58));
\GRLFPC20_COMB_V_E_STDATA_1_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(3),
dataa => \GRLFPC20.R.FSR.CEXC\(3),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(35));
\GRLFPC20_COMB_V_E_STDATA_1_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(14),
dataa => \GRLFPC20.R.FSR.FTT\(0),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(46));
\GRLFPC20_COMB_V_E_STDATA_1_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(11),
dataa => CPO_CCZ(1),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(47),
datac => \GRLFPC20.FPI.OP2_X\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(45),
datac => \GRLFPC20.FPI.OP2_X\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(44),
datac => \GRLFPC20.FPI.OP2_X\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(41),
datac => \GRLFPC20.FPI.OP2_X\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(174),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2_REP1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(53),
datac => \GRLFPC20.FPI.OP2_X\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(51),
datac => \GRLFPC20.FPI.OP2_X\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(0),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(40),
dataa => N_702,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(156),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(42),
dataa => N_700,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(158),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(44),
dataa => N_698,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(160),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(48),
dataa => N_694,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(164),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(50),
dataa => N_692,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(166),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(53),
datac => \GRLFPC20.FPI.OP1_X\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(63),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(52),
datac => \GRLFPC20.FPI.OP1_X\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(66),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(49),
datac => \GRLFPC20.FPI.OP1_X\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(73),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(42),
datac => \GRLFPC20.FPI.OP1_X\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(76),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(39),
datac => \GRLFPC20.FPI.OP1_X\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(79),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(36),
datac => \GRLFPC20.FPI.OP1_X\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(80),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(35),
datac => \GRLFPC20.FPI.OP1_X\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(251),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(61),
datac => \GRLFPC20.FPI.OP1_X\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(256),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(53),
datac => \GRLFPC20.FPI.OP1_X\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(257),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(52),
datac => \GRLFPC20.FPI.OP1_X\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(27));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(22));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111111010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_SLCONTROL_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111111100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_1\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(49),
dataa => N_693,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(165),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(51),
dataa => N_691,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(167),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(69),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(46),
datac => \GRLFPC20.FPI.OP1_X\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(72),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(43),
datac => \GRLFPC20.FPI.OP1_X\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(40),
datac => \GRLFPC20.FPI.OP1_X\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(78),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(37),
datac => \GRLFPC20.FPI.OP1_X\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(19));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111001100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_A_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20_A\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SRCONTROL_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(254),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(58),
datac => \GRLFPC20.FPI.OP1_X\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(26),
dataa => N_716,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(28),
dataa => N_714,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(144),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(33),
dataa => N_709,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(149),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(34),
dataa => N_708,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(150),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(37),
dataa => N_705,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(153),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(38),
dataa => N_704,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(154),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(39),
dataa => N_703,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(155),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(41),
dataa => N_701,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(157),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(52),
datac => \GRLFPC20.FPI.OP2_X\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(49),
datac => \GRLFPC20.FPI.OP2_X\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(46),
datac => \GRLFPC20.FPI.OP2_X\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(43),
datac => \GRLFPC20.FPI.OP2_X\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(40),
datac => \GRLFPC20.FPI.OP2_X\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(38),
datac => \GRLFPC20.FPI.OP2_X\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(37),
datac => \GRLFPC20.FPI.OP2_X\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(35),
datac => \GRLFPC20.FPI.OP2_X\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(372),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(27),
dataa => N_715,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(143),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(32),
dataa => N_710,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(148),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(36),
dataa => N_706,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(152),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(47),
dataa => N_695,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(163),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(52),
dataa => N_690,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(168),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(48),
datac => \GRLFPC20.FPI.OP2_X\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(39),
datac => \GRLFPC20.FPI.OP2_X\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(36),
datac => \GRLFPC20.FPI.OP2_X\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(45),
dataa => N_697,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(161),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(62));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_35\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_56\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_56\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_18\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_55\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_55\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_54\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_54\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_50\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_50\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_48\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(46));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100100111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_45\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_30\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_43\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_43\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_43\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_42\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_41\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_35\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_34\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_34\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_32\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_31\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_30\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_28\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_28\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0_62__ROM\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_27\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_24\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_24\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_12\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_12\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_15\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_18\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_14\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_14\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_14\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_14\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_13\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_11\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_11\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_11\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_9\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_7\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_7\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0_62__ROM\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0_62__ROM\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(62));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_58\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_57\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_57\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_57\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_56\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_56\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_56\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_56\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_55\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_55\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_55\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_54\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_54\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_54\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_53\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_50\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_50\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_49\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_13\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_48\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_43\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_42\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_42\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(40));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100100111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_36\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_35\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_34\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_34\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_33\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_31\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_31\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_30\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_58\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_28\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_27\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_22\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110010000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_15\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_14\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_14\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_14\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_13\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_11\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_9\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_7\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(61),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_60\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(60),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_59\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_59\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_57\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_57\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_55\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_55\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_55\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_50\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_50\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_50\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_49\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_48\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_48\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_43\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_43\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_42\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_42\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_16\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_37\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_34\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_34\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_33\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_31\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_31\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_30\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011000110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_27\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_27\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011000110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110010000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_13\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_13\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_10\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_7\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_7\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_0\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110010000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_61\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(62));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_58\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_57\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_56\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_55\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011110100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_55\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100100111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_54\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_20\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_50\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_50\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_48\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_48\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_44\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(44));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011000110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_43\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_42\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(43));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_42\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_42\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_37\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_34\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_34\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_34\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_33\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_31\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_30\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_30\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(30));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_29\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_28\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(29));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_28\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_27\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_27\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_26\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_26\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_25\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_22\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(23));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_19\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_14\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(15));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_14\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_14\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(11));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_9\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_9\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_8\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_16\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011000110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_7\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(7));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_6\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_5\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_4\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(4));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_3\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_1\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110001001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000011011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011001010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0_62__ROM\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\);
\GRLFPC20_R_E_STDATA_RNO_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_0__G2\,
dataa => \GRLFPC20.R.FSR.CEXC\(0),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(32));
\GRLFPC20_R_E_STDATA_RNO_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_1__G2\,
dataa => \GRLFPC20.R.FSR.CEXC\(1),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(33));
\GRLFPC20_R_E_STDATA_RNO_0_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110011111010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_17__G2\,
dataa => N_609,
datab => N_673,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_R_E_STDATA_RNO_0_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_20__G2\,
dataa => N_612,
datab => N_676,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_R_E_STDATA_RNO_0_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_21__G2\,
dataa => N_613,
datab => N_677,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_R_E_STDATA_RNO_0_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_29__G2\,
dataa => N_621,
datab => N_685,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_21_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101101000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_21\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(42),
datac => \GRLFPC20.FPI.OP2_X\(39));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(273),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(60),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(60));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110100001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(258),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(259),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(111),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(111));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_SELECTQUOBITS_QUOBITS_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000111100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.QUOBITS\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111111010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(21));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(110),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(110));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(108),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(108));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(95),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(95));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(70),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(45),
datac => \GRLFPC20.FPI.OP1_X\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(67),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(48),
datac => \GRLFPC20.FPI.OP1_X\(45));
\GRLFPC20_COMB_V_E_STDATA_1_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(16),
dataa => \GRLFPC20.R.FSR.FTT\(2),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(48));
GRLFPC20_COMB_V_I_V_1_F1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111111110100")
port map (
combout => \GRLFPC20.COMB.V.I.V_1_F1\,
dataa => N_3,
datab => \GRLFPC20.R.I.V\,
datac => \GRLFPC20.COMB.UN2_HOLDN\,
datad => \GRLFPC20.COMB.UN19_IUEXEC\);
\GRLFPC20_COMB_RS1_1_0_X_RNI5ER71_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100000001000")
port map (
combout => \GRLFPC20.COMB.V.A.RF1REN_1_670_I_M4\,
dataa => N_68,
datab => \GRLFPC20.RS1V_0_SQMUXA\,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.COMB.RS1_1_0_X\(0));
\GRLFPC20_COMB_RS1_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110000000")
port map (
combout => \GRLFPC20.COMB.RS1_1\(0),
dataa => N_68,
datab => \GRLFPC20.RS1V_0_SQMUXA\,
datac => \GRLFPC20.COMB.RS1_1_SN_M2_X\,
datad => \GRLFPC20.COMB.RS1_1_0_X\(0));
\GRLFPC20_COMB_RS1_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110000000")
port map (
combout => \GRLFPC20.COMB.RS1_1\(2),
dataa => N_70,
datab => \GRLFPC20.RS1V_0_SQMUXA\,
datac => \GRLFPC20.COMB.RS1_1_SN_M2_X\,
datad => \GRLFPC20.COMB.RS1_1_0_X\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(30),
dataa => N_712,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(146),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(314),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(311),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(256),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(256));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(253),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(59),
datac => \GRLFPC20.FPI.OP1_X\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(250),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(62),
datac => \GRLFPC20.FPI.OP1_X\(59));
\GRLFPC20_COMB_V_E_STDATA_1_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(30),
dataa => \GRLFPC20.R.FSR.RD\(0),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(62));
\GRLFPC20_COMB_V_E_STDATA_1_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(27),
dataa => \GRLFPC20.R.FSR.TEM\(4),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(59));
\GRLFPC20_COMB_DBGDATA_4_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(19),
dataa => N_611,
datab => N_675,
datac => N_391,
datad => N_390);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010111010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_I_0_0__G0_0_M2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_RNO_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101010100010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SCTRL_NEW_0_0__G0_I_M2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SRCONTROL_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SRCONTROL_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SRCONTROL_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100010011000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(13));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SRONEMORE: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRONEMORE\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(2),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(255),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(255));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(254),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(254));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_249_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(249),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(249));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(252),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(252));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(250),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(250));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(50),
datac => \GRLFPC20.FPI.OP2_X\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(265),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111111010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(8));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101111111010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(313),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(267),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_R_E_STDATA_RNO_0_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_19__G2\,
dataa => N_611,
datab => N_675,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(31),
dataa => N_711,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(147),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(255),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(57),
datac => \GRLFPC20.FPI.OP1_X\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(64),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(51),
datac => \GRLFPC20.FPI.OP1_X\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(61),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(51),
datac => \GRLFPC20.FPI.OP1_X\(54));
\GRLFPC20_COMB_V_E_STDATA_1_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(25),
dataa => \GRLFPC20.R.FSR.TEM\(2),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(57));
\GRLFPC20_COMB_V_E_STDATA_1_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(22),
dataa => \GRLFPC20.R.FSR.NONSTD\,
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(32));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(91),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(91));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(43),
dataa => N_699,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(159),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP1\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(16));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(102),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(102));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(101),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(101));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(278),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(299),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(301),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_RNDMODESELECT_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110011101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
datab => \GRLFPC20.FPI.LDOP\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(77),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(38),
datac => \GRLFPC20.FPI.OP1_X\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(74),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(41),
datac => \GRLFPC20.FPI.OP1_X\(38));
\GRLFPC20_COMB_V_E_STDATA_1_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(9),
dataa => \GRLFPC20.R.FSR.AEXC\(4),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(41));
\GRLFPC20_COMB_V_E_STDATA_1_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(6),
dataa => \GRLFPC20.R.FSR.AEXC\(1),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(38));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(251),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(251));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_12_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_12\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49));
\GRLFPC20_COMB_V_E_STDATA_1_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(31),
dataa => \GRLFPC20.R.FSR.RD\(1),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(63));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_245_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(245),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
datab => NN_1,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(53),
dataa => N_689,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(169),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_25_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_25\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_WAITMULXFF_UN2_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010011110100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.UN2_TEMP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(46),
dataa => N_696,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(162),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_NOTABORTNULLEXC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000111110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.NOTABORTNULLEXC\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_246_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(246),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(246));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_247_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(247),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(247));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M2_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111011111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M2_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M5_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M5_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M8_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M8_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M11_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001000110010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M11_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110011011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(54),
dataa => N_688,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(170),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(24));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(49));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111010111110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M11_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M11\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPYBUS_2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_S_8_20_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110111111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_S_8_20\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_REP2\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIGKP11_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110100001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL_SN_M3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(240),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(59),
datac => \GRLFPC20.FPI.OP2_X\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(241),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(58),
datac => \GRLFPC20.FPI.OP2_X\(55));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(242),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(57),
datac => \GRLFPC20.FPI.OP2_X\(54));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(238),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(61),
datac => \GRLFPC20.FPI.OP2_X\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(3),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_248_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(248),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(248));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(244),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(55),
datac => \GRLFPC20.FPI.OP2_X\(52));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(257),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(257));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_SFTLFT_UN4_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100011111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.UN4_TEMP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010100110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(243),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(56),
datac => \GRLFPC20.FPI.OP2_X\(53));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(239),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(60),
datac => \GRLFPC20.FPI.OP2_X\(57));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_33_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_33\(237),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(62),
datac => \GRLFPC20.FPI.OP2_X\(59));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(5));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_2\(253),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(253));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(20));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(277),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_COMB_DBGDATA_4_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(28),
dataa => N_620,
datab => N_684,
datac => N_391,
datad => N_390);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_41_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_41\(252),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(60),
datac => \GRLFPC20.FPI.OP1_X\(57));
\GRLFPC20_R_E_STDATA_RNO_0_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_28__G2\,
dataa => N_620,
datab => N_684,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIRVP11_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STATUS\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39));
\GRLFPC20_R_I_CC_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011100000")
port map (
combout => \GRLFPC20.R.I.CC_0_0_0__G4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38));
\GRLFPC20_R_I_CC_RNO_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010110000")
port map (
combout => \GRLFPC20.R.I.CC_0_0_1__G4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38));
\GRLFPC20_COMB_RS2_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011001110000000")
port map (
combout => \GRLFPC20.COMB.RS2_1\(0),
dataa => N_43,
datab => N_3,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.R.A.RS2\(0));
\GRLFPC20_COMB_RS2_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011001110000000")
port map (
combout => \GRLFPC20.COMB.RS2_1\(2),
dataa => N_45,
datab => N_3,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.R.A.RS2\(2));
GRLFPC20_COMB_FPDECODE_ST3_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.COMB.FPDECODE.ST3_1\,
dataa => N_65,
datab => N_66,
datac => N_64,
datad => N_67);
\GRLFPC20_COMB_DBGDATA_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011100100")
port map (
combout => CPO_DBG_DATAZ(13),
dataa => N_390,
datab => \GRLFPC20.COMB.DBGDATA_4_0_X\(13),
datac => \GRLFPC20.R.STATE\(1),
datad => \GRLFPC20.R.STATE\(0));
\GRLFPC20_COMB_V_E_STDATA_1_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111100100000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(13),
dataa => \GRLFPC20.R.STATE\(1),
datab => \GRLFPC20.R.STATE\(0),
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.FPI.OP1_X\(45));
\GRLFPC20_COMB_RS2_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011001110000000")
port map (
combout => \GRLFPC20.COMB.RS2_1\(3),
dataa => N_46,
datab => N_3,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.R.A.RS2\(3));
\GRLFPC20_R_E_STDATA_RNO_0_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111110011111010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_18__G2\,
dataa => N_610,
datab => N_674,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_R_E_STDATA_RNO_0_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110000001010")
port map (
combout => \GRLFPC20.R.E.STDATA_1_0_12__G2\,
dataa => N_604,
datab => N_668,
datac => \GRLFPC20.R.A.AFSR\,
datad => \GRLFPC20.COMB.UN1_R.A.RS1_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(71),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(44),
datac => \GRLFPC20.FPI.OP1_X\(41));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(68),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(44),
datac => \GRLFPC20.FPI.OP1_X\(47));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_19_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(65),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP1_X\(50),
datac => \GRLFPC20.FPI.OP1_X\(47));
\GRLFPC20_COMB_V_E_STDATA_1_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.COMB.V.E.STDATA_1_1\(15),
dataa => \GRLFPC20.R.FSR.FTT\(1),
datab => \GRLFPC20.R.A.AFSR\,
datac => \GRLFPC20.FPI.OP1_X\(47));
\GRLFPC20_COMB_DBGDATA_4_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(12),
dataa => N_604,
datab => N_668,
datac => N_391,
datad => N_390);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_A_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100100111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_A\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_36\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_36\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(37));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_6_A_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_6_A\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_36\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_36\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_A_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011000110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10_A\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_17\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_17\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110010000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_10_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_10\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(18));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_17\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000100100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_17\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_13_A_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001101100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_13_A\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_31\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_35\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_S_CMP_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.S_CMP_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81));
\GRLFPC20_R_I_EXC_RNO_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100001010")
port map (
combout => \GRLFPC20.R.I.EXC_2_0_5__G0\,
dataa => \GRLFPC20.R.I.EXC\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(69),
datac => \GRLFPC20.COMB.UN2_HOLDN\,
datad => \GRLFPC20.COMB.UN19_IUEXEC\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(53));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN25_NOTXZYFROMD: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(12));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN8_TEMP_2_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100011110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_2\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_2_A\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN8_TEMP_2_A_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010111110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN8_TEMP_2_A\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(35),
dataa => N_707,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(151),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(48));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(26));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(45));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(200),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_SN_M2\,
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(35));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(34));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(93),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(93));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(85),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(83),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(83));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(293),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_COMB_RS2_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011001110000000")
port map (
combout => \GRLFPC20.COMB.RS2_1\(1),
dataa => N_44,
datab => N_3,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.R.A.RS2\(1));
\GRLFPC20_COMB_RS1_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110000000")
port map (
combout => \GRLFPC20.COMB.RS1_1\(4),
dataa => N_72,
datab => \GRLFPC20.RS1V_0_SQMUXA\,
datac => \GRLFPC20.COMB.RS1_1_SN_M2_X\,
datad => \GRLFPC20.COMB.RS1_1_0_X\(4));
\GRLFPC20_COMB_RS1_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000111110000000")
port map (
combout => \GRLFPC20.COMB.RS1_1\(3),
dataa => N_71,
datab => \GRLFPC20.RS1V_0_SQMUXA\,
datac => \GRLFPC20.COMB.RS1_1_SN_M2_X\,
datad => \GRLFPC20.COMB.RS1_1_0_X\(3));
\GRLFPC20_COMB_RS2_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011001110000000")
port map (
combout => \GRLFPC20.COMB.RS2_1\(4),
dataa => N_47,
datab => N_3,
datac => \GRLFPC20.RS2_0_SQMUXA\,
datad => \GRLFPC20.R.A.RS2\(4));
\GRLFPC20_COMB_DBGDATA_4_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011001010")
port map (
combout => CPO_DBG_DATAZ(20),
dataa => N_612,
datab => N_676,
datac => N_391,
datad => N_390);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_3_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101011001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_3\(29),
dataa => N_713,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(145),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datad => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_4_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(28));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_DPATH_NEW_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_1\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
datab => \GRLFPC20.FPI.OP2_X\(54),
datac => \GRLFPC20.FPI.OP2_X\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M2_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2\(87),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M2S2_REP1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(87));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(283),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(287),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_SN_M1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_115_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(115),
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_DPATH_NEW_7_SQMUXA_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_NEW_7_SQMUXA_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_32_0_RNIPG1G_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_M1_0_A2_0_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_ENTRYSHFT_UN3_S_SQRT_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN3_S_SQRT_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNIVRM8_221_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(221),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_RNI40M8_217_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_E_3_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(217),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_INEXACTSIG_UN13_INEXACT_10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.INEXACTSIG.UN13_INEXACT_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_SELINITREMBIT_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELINITREMBIT_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN4_NOTSHIFTCOUNT1_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN4_NOTSHIFTCOUNT1_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(14));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_31_S_0_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31_S_0\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_AEBEEXC_UN3_NOTAZERODENORM_0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.AEBEEXC.UN3_NOTAZERODENORM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN25_NOTXZYFROMD_RNIIJIB1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M2_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_M1_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_2_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_3_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL_I_M_0\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_PCTRL_NEW_43_2_C\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_32_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_32_0\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_31\(75));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_PCTRL_NEW_12_30_S_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_12_30_S\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50));
GRLFPC20_R_MK_HOLDN2_RNILNJ1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => CPO_HOLDNZ,
dataa => \GRLFPC20.R.MK.HOLDN2\,
datab => \GRLFPC20.R.MK.HOLDN1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(362),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(359),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(358),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(356),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(354),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(349),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(345),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(341),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(333),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(332),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(331),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(330),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(327),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(323),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(322),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(321),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_I_O2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_I_O2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_ROMXZSL2FROMC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.ROMXZSL2FROMC\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_3_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_3_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(1));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_UN38_SHDVAR_3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.UN38_SHDVAR_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIP4QM_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.ENTRYSHFT.UN6_S_0_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(61),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(63),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(64),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(65),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(66),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(67),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(68),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(69),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(70),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(71),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(72),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(73),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(74),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(76),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(77),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(78),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(79),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(80),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(81),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(82),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(84),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(86),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(88),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(89),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(90),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(92),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(94),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(96),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(97),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(98),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(99),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(100),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(103),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(104),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(105),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(106),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(107),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(109),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(112),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_61_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(61),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_63_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(63),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_64_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(64),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_65_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(65),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_66_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(66),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_67_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(67),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_68_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(68),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(69),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_70_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(70),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_71_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(71),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_72_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(72),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_73_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(73),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(74),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_75_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(75),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_76_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(76),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_77_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(77),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_78_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(78),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_79_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(79),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(80),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_81_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(81),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_82_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(82),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_84_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(84),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_86_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(86),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_88_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(88),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_89_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(89),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_90_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(90),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_92_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(92),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_94_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(94),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_96_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(96),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_97_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(97),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_98_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(98),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_99_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(99),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_100_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(100),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_103_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(103),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_104_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(104),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_105_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(105),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_106_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(106),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_107_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(107),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_109_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(109),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_112_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(112),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_115_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(115),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_SUB_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000111010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SUB\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(18),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(46),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_118_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_118\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_125_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_125\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_2_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(16),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_134_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_134\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_12_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_12\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_12_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_12\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_11_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_49\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_11_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_57\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_11_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_11_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_31\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_31\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_11_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_11\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_9_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_61\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_38\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_9_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_43\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_9_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_15\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_9_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_9_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_53\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_48\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_48\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_46\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(40),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_32\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_19\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_31\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_27\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_27\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_8_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_8\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_62_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(62),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_61\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_61\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_38\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_37\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_37\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_9\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_9\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_5_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_5\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_4_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_49\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_4_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_54\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_20\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_4_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_44\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_49\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_4_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(15),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_14\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_14\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_4_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_4_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_4_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_4\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_57\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_35\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_33\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_16\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_2_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_2\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_47\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_58\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_1_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_56\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_1_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_1\(11),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_10\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_EXPBREGLOADEN_RNIG92H: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3\,
dataa => \GRLFPC20.FPI.LDOP\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIVU6R_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
datab => \GRLFPC20.FPI.LDOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(41),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(60),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_60_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(60),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(57),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_113_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(113),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(111),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_113_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(113),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_111_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(111),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_T_3_RNO_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.NOTDIVC\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLCREGXZ_UN1_INFORCREGDB: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLCREGXZ.UN1_INFORCREGDB\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(17),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(110),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(108),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(95),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_110_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(110),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_108_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(108),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_95_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(95),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(54),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(319),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(18),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(355),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(365),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(22),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(351),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(352),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(353),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(369),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_256_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(256),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_58_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(58),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_XZXBUS_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(43),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_TEMP: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TEMP\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_255_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(255),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_254_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(254),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_249_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(249),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD9\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_252_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(252),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_250_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(250),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_59_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(59),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(14),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(19),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(21),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(51),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(52),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110111011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(2),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(2));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(29),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(344),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(30),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(343),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(342),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(337),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(373),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_114_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(114),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(367),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(32),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(91),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_91_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(91),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(56),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(317),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(320),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(47),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(326),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(44),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(329),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(39),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(334),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(38),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(335),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(37),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(336),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(27),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(346),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(347),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(25),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(348),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(23),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(350),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(13),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(360),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(361),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_0_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101110001011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5_0\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(312),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_DPATH_0_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.DPATH_0\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(12),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(50),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(42),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(102),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(101),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_102_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(102),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_101_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(101),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIRPTN_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIQOTN_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_251_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(251),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_74_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_18_0_74__G0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(62),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => NN_1,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_SELECTQUOBITS_NOTDIVC_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.SELECTQUOBITS.NOTDIVC\(1),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110110001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(55),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(339),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(33),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(340),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_246_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(246),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_247_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(247),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD11\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M5S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M5S2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_COUNTSUCCESSIVEZERO_M8S2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.COUNTSUCCESSIVEZERO_M8S2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_COMPUTECONST_UN25_RESVEC_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.COMPUTECONST.UN25_RESVEC_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(24),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_LEFTSHIFTERBL_S_8_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.S_8\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_2_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_2_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_2_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPXBUS_2_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_2\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_EXPYBUS_0_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.EXPYBUS_0\(4),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_EXPYBUS_2_1_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2_1\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_GRFPUELOC_0_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC_0\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.SLCONTROL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNILV5N1_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_0_I\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_240_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(240),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD4\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_241_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(241),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_242_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(242),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_235_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(235),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD9\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_238_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(238),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD6\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(3),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_248_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(248),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_244_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(244),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_257_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(257),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_TOPBITSIN_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.TOPBITSIN\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_236_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(236),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD8\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_234_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(234),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD10\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_232_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(232),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(5),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_253_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(253),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_243_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(243),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_239_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(239),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD5\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_237_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1\(237),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD7\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_0_232_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0\(232),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPAREGLOADEN_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_SFTLFT_AREGXORBREG: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.AREGXORBREG\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_SXC_SFTLFT_UN1_GRFPUS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SFTLFT.UN1_GRFPUS\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(24));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_PXS_FEEDBACKMULXFF_UN7_FEEDBACK_1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.FEEDBACKMULXFF.UN7_FEEDBACK_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(20),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD3\);
GRLFPC20_FPI_LDOP_2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.FPI.LDOP_2\,
dataa => \GRLFPC20.R.MK.RST2\,
datab => \GRLFPC20.R.MK.RST\);
GRLFPC20_COMB_LOCKGEN_DEPCHECK_RNO: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100010001")
port map (
combout => \GRLFPC20.ANNULRES_0_SQMUXA_12_1\,
dataa => \GRLFPC20.R.I.EXEC\,
datab => \GRLFPC20.R.E.FPOP\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIGJHM_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STATUS\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DECODESTATUS_UN7_STATUS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DECODESTATUS.UN7_STATUS\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38));
GRLFPC20_COMB_QNE2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => \GRLFPC20.COMB.QNE2\,
dataa => \GRLFPC20.R.STATE\(0),
datab => \GRLFPC20.R.STATE\(1));
GRLFPC20_COMB_PEXC12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000100")
port map (
combout => CPO_EXCZ,
dataa => \GRLFPC20.R.STATE\(1),
datab => \GRLFPC20.R.STATE\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNO_0_69_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G0_I_O4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_MUX_9_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110010011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_9\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_35\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RNIHTQM_80_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011001100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.ENTRYSHFT.S_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81));
GRLFPC20_COMB_UN19_IUEXEC_RNIIF5I: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.G_884\,
dataa => \GRLFPC20.COMB.UN2_HOLDN\,
datab => \GRLFPC20.COMB.UN19_IUEXEC\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(53),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_UN26_XZYBUSLSBS: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN26_XZYBUSLSBS\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(231),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN25_NOTXZYFROMD\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN15_XZROUNDOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN15_XZROUNDOUT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_UN23_XZROUNDOUT: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110111011101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN23_XZROUNDOUT\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_EXPADDERSHFT_MIXOIN_0_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.MIXOIN\(0),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(26),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_FAX_TEMP_1_0_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_1_0\(31),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN3_NOTXZYFROMD\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_RIGHTSHIFTERBL_S_8_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001101010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.RIGHTSHIFTERBL.S_8\(6),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SRCONTROL_1\(3));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(35),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(34),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(93),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(85),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(83),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_93_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(93),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_85_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(85),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_83_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(83),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_1_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100011011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_1\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(36),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_1_2_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110001011100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_2\(28),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD3\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M1_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010110010101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M1\(87),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.DPATH_M2\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_RIN_DPATH_M0_87_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100101011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M0\(87),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\,
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZBREGLOADEN_REP1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(49),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(48),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(325),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(45),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(328),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(10),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(363),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_MIXOIN_3_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.MIXOIN_3\(9),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(364),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0));
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100101101001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_11\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD11\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_10\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD10\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_9\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD9\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_8\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD8\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_7\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD7\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_6\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD6\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_5\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD5\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_4\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD4\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD3\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_GRFPUE_ADD0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.GRFPUE_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
cin => N_19200);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(8),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
datab => GND,
cin => N_10425);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110110001101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(7),
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
cin => N_10424);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(6),
cout => N_10425,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
cin => N_10423);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_5_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110110010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(5),
cout => N_10424,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
cin => N_10422);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_4_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(4),
cout => N_10423,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
cin => N_10421);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_3_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110110010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(3),
cout => N_10422,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
cin => N_10419);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_2_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0101101010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(2),
cout => N_10421,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
cin => N_10418);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_A_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0000000000100010")
port map (
cout => N_10418,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN1_R_PCTRL_1_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001100100100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.PCTRL\(1),
cout => N_10419,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.WAITMULXFF.NOTSAMPLEDWAIT\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD57: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100101101001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(57),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(57),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_56\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD56: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(56),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(56),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_55\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD55: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(55),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(55),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_54\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD54: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(54),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(54),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_53\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD53: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_53\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(53),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(53),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_52\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD52: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_52\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(52),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(52),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_51\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD51: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_51\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(51),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(51),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_50\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD50: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(50),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(50),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_49\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD49: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_49\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(49),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(49),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_48\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD48: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(48),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(48),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_47\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD47: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_47\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(47),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(47),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_46\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD46: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_46\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(46),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(46),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_45\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD45: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_45\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(45),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(45),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_44\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD44: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(44),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(44),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_43\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD43: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(43),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(43),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_42\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD42: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(42),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(42),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_41\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD41: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_41\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(41),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(41),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_40\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD40: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_40\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(40),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(40),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_39\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD39: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_39\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(39),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(39),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_38\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD38: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_38\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(38),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(38),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_37\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD37: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_37\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(37),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(37),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_36\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD36: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(36),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(36),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_35\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD35: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_35\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(35),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(35),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_34\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD34: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(34),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(34),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_33\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD33: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_33\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(33),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(33),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_32\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD32: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_32\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(32),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(32),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_31\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD31: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_31\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(31),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(31),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_30\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD30: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(30),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(30),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_29\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD29: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(29),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(29),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_28\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD28: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(28),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(28),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_27\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD27: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(27),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(27),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_26\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD26: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_26\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(26),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(26),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_25\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD25: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(25),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(25),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_24\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_24\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(24),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(24),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_23\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD23: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_23\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(23),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(23),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_22\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD22: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(22),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(22),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_21\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD21: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_21\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(21),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(21),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_20\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD20: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_20\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(20),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(20),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_19\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD19: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_19\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(19),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(19),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_18\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD18: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_18\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(18),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(18),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_17\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD17: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_17\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(17),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(17),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_16\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD16: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_16\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(16),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(16),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_15\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_15\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(15),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(15),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_14\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(14),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(14),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_13\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD13: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(13),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(13),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_12\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(12),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_11\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(11),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_10\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(10),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_9\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(9),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_8\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(8),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_7\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(7),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_6\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(6),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_5\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(5),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_4\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(4),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUF_ADD0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "0110100111010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.TEMP_2\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.XZXBUS\(0),
cin => N_19201);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011010010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(12),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(12),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_11\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD11: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD11\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(11),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(11),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_10\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD10: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD10\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(10),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(10),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_9\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD9\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(9),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(9),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_8\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD8\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(8),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(8),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_7\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD7\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(7),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(7),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_6\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD6: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD6\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(6),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(6),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_5\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD5\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(5),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(5),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_4\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD4\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(4),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(4),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_3\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD3\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(3),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(2),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(1),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_0\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_UN6_GRFPUE_ADD0: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPXBUS_3\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.GRFPUELOC_0\(0),
cin => N_19202);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_1_RNIOH979: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD3\,
cout => N_19203,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_1_RNI4VBC4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_2_RNI1UBL1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFI1H_51_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(51),
cin => N_19204);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_2_RNI92KV9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD3\,
cout => N_19205,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_RNI4EUH4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_1_RNIFOE02: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI2BTI_52_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(52),
cin => N_19206);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_47_TRFWWBASICCELL_TEMP2_3_RNICTUGA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD3\,
cout => N_19207,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_2_RNIJOO15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_2_RNIGJJS1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNITL6P_53_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(53),
cin => N_19208);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_48_TRFWWBASICCELL_TEMP2_3_RNIOAK3A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD3\,
cout => N_19209,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_RNI5IB05: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_1_RNICEO82: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI1F4S_54_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(54),
cin => N_19210);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_49_TRFWWBASICCELL_TEMP2_3_RNI067S8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD3\,
cout => N_19211,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_3_RNIUEGH4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_1_RNIINH12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI282V_55_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(55),
cin => N_19212);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_50_TRFWWBASICCELL_TEMP2_RNIIMEO9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD3\,
cout => N_19213,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_2_RNICM064: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_2_RNIR0BQ1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI610I_56_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(56),
cin => N_19214);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_51_TRFWWBASICCELL_TEMP2_RNIMIFAC: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD3\,
cout => N_19215,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.SI_118_1.SUM\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_52_TRFWWBASICCELL_TEMP2_3_RNIA8195: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_61_1.SUM_0_A2\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_53_TRFWWBASICCELL_TEMP2_3_RNI084J1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.CI_2_SUM0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9QTK_57_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(57),
cin => N_19216);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_2_RNI90IR7: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD3\,
cout => N_19217,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_1_RNIF7DS3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_1_RNID06M1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI19IG_36_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(36),
cin => N_19218);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_3_RNI86OH8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD3\,
cout => N_19219,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_RNIFVEL3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_2_RNIK9VE1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI32GJ_37_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(37),
cin => N_19220);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_32_TRFWWBASICCELL_TEMP2_3_RNIV0AK9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD3\,
cout => N_19221,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_RNICMLF4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_3_RNISION1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI6RDM_38_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(38),
cin => N_19222);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_33_TRFWWBASICCELL_TEMP2_1_RNI5SV2A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD3\,
cout => N_19223,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_RNI533L4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_3_RNIGBJ02: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9KBP_39_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(39),
cin => N_19224);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_34_TRFWWBASICCELL_TEMP2_1_RNIOP1MA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD3\,
cout => N_19225,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_RNIJQDB5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_RNIKAJ42: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIPSAS_40_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(40),
cin => N_19226);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_35_TRFWWBASICCELL_TEMP2_1_RNIOGM2A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD3\,
cout => N_19227,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_1_RNIN9755: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_3_RNITDBE2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIUL8V_41_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(41),
cin => N_19228);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_36_TRFWWBASICCELL_TEMP2_3_RNI4RA0A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD3\,
cout => N_19229,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_RNIIQ4L4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_RNI7BV02: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFFAU_42_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(42),
cin => N_19230);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_37_TRFWWBASICCELL_TEMP2_2_RNIMAHU9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD3\,
cout => N_19231,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_2_RNI0TTV4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_3_RNI73HQ1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIPPFO_43_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(43),
cin => N_19232);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_38_TRFWWBASICCELL_TEMP2_1_RNI4MR69: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD3\,
cout => N_19233,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_1_RNI4JDG4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_RNI3RK92: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNISIDR_44_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(44),
cin => N_19234);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_39_TRFWWBASICCELL_TEMP2_2_RNI2QIA8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD3\,
cout => N_19235,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_2_RNIEHA54: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_RNIB23O1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFOFT_45_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(45),
cin => N_19236);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_40_TRFWWBASICCELL_TEMP2_3_RNITQ8H8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD3\,
cout => N_19237,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_2_RNI00714: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_1_RNIKG8O1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI359H_46_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(46),
cin => N_19238);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_41_TRFWWBASICCELL_TEMP2_3_RNIPU129: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD3\,
cout => N_19239,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_2_RNIG9N54: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_1_RNISP1H1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI7U6K_47_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(47),
cin => N_19240);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_42_TRFWWBASICCELL_TEMP2_3_RNIC4DV9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD3\,
cout => N_19241,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_RNIRC2F4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_1_RNI33RP1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIAN4N_48_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(48),
cin => N_19242);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_43_TRFWWBASICCELL_TEMP2_3_RNIVTLE9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD3\,
cout => N_19243,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_RNI2O405: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_2_RNINRL22: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIDG2Q_49_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(49),
cin => N_19244);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_44_TRFWWBASICCELL_TEMP2_2_RNI1SQT8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD3\,
cout => N_19245,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_45_TRFWWBASICCELL_TEMP2_RNIDFDB4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_46_TRFWWBASICCELL_TEMP2_RNI9PA22: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNISO1T_50_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(50),
cin => N_19246);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_2_RNIS4ES9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD3\,
cout => N_19247,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_RNI7F125: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_1_RNIRN962: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI644V_21_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(21),
cin => N_19248);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_3_RNIS09P9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD3\,
cout => N_19249,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_2_RNI7PBJ4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_2_RNIBC512: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI9RMN_22_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(22),
cin => N_19250);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_17_TRFWWBASICCELL_TEMP2_RNI0404A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD3\,
cout => N_19251,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_3_RNI5KUR4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_2_RNI9LLQ1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIK12N_23_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(23),
cin => N_19252);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_18_TRFWWBASICCELL_TEMP2_1_RNIDGMNA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD3\,
cout => N_19253,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_3_RNISSGV4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_1_RNI7GQ62: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI6D9U_24_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(24),
cin => N_19254);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_19_TRFWWBASICCELL_TEMP2_1_RNIV0RCA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD3\,
cout => N_19255,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_3_RNI1IB85: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_1_RNIV6AB2: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIRJTS_25_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(25),
cin => N_19256);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_20_TRFWWBASICCELL_TEMP2_RNIKVCQ9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD3\,
cout => N_19257,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_2_RNIDMN15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_1_RNIKSB92: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNITCRV_26_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(26),
cin => N_19258);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_21_TRFWWBASICCELL_TEMP2_3_RNI7TJD9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD3\,
cout => N_19259,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_2_RNIEJVG4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_RNIBKO12: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFI1O_27_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(27),
cin => N_19260);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_22_TRFWWBASICCELL_TEMP2_RNISAPE9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD3\,
cout => N_19261,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_3_RNIDHLG4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_3_RNIK2ML1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3VML_28_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(28),
cin => N_19262);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_23_TRFWWBASICCELL_TEMP2_1_RNIIIT0A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD3\,
cout => N_19263,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_1_RNIKP8L4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_3_RNI8RGU1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI5OKO_29_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(29),
cin => N_19264);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_24_TRFWWBASICCELL_TEMP2_2_RNITT8G9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD3\,
cout => N_19265,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_1_RNIIIQP4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_2_RNISJB72: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIM0KR_30_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(30),
cin => N_19266);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_25_TRFWWBASICCELL_TEMP2_RNIK7719: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD3\,
cout => N_19267,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_3_RNITDMH4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_3_RNI5T402: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIPPHU_31_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(31),
cin => N_19268);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_26_TRFWWBASICCELL_TEMP2_RNIBDC59: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD3\,
cout => N_19269,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_2_RNIPQTC4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_2_RNI4O9S1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNITIFH_32_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(32),
cin => N_19270);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_27_TRFWWBASICCELL_TEMP2_RNIED6P8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD3\,
cout => N_19271,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_RNIJU8D4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_1_RNI1JEO1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIOTON_33_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(33),
cin => N_19272);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_28_TRFWWBASICCELL_TEMP2_3_RNIUDDV8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD3\,
cout => N_19273,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_3_RNIR5584: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_RNIE0RT1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIQMMQ_34_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(34),
cin => N_19274);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_29_TRFWWBASICCELL_TEMP2_RNI19488: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD3\,
cout => N_19275,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_30_TRFWWBASICCELL_TEMP2_1_RNIGEP64: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_31_TRFWWBASICCELL_TEMP2_RNIM79S1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNITFKT_35_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(35),
cin => N_19276);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_0_TRFWWBASICCELL_TEMP2_2_RNIHPCSA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD3\,
cout => N_19277,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.REMWTAGE57.0.TRFWWBASICCELL.CIN_4\,
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_1_RNI4K1C5: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_1_RNIN5G82: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIMA741_6_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(6),
cin => N_19278);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_1_TRFWWBASICCELL_TEMP2_3_RNIS0B5A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD3\,
cout => N_19279,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_2_RNILNG15: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_3_RNIIS472: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIBH0T_7_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(7),
cin => N_19280);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_2_TRFWWBASICCELL_TEMP2_RNIV6LT8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD3\,
cout => N_19281,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_1_RNID42I4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_1\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI6I1B2_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIEAUV_8_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(8),
cin => N_19282);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_3_TRFWWBASICCELL_TEMP2_2_RNIBESB8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD3\,
cout => N_19283,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_1_RNI9ID24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_RNIAIOK1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIVFVT_9_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(9),
cin => N_19284);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_4_TRFWWBASICCELL_TEMP2_RNIIBQE8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD3\,
cout => N_19285,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_1_RNI79R14: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_2_RNI19FO1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI259H_10_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(10),
cin => N_19286);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_5_TRFWWBASICCELL_TEMP2_2_RNIR4PF8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD3\,
cout => N_19287,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_3_RNI08K24: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_2_RNI7I8H1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI4U6K_11_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(11),
cin => N_19288);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_6_TRFWWBASICCELL_TEMP2_1_RNI6C739: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD3\,
cout => N_19289,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_1_RNIURLV3: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_3_RNINGAM1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI7N4N_12_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(12),
cin => N_19290);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_7_TRFWWBASICCELL_TEMP2_RNIMGO99: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD3\,
cout => N_19291,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_RNIBO4J4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_3_RNI6FCR1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNII5BM_13_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(13),
cin => N_19292);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_8_TRFWWBASICCELL_TEMP2_1_RNIB5F09: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD3\,
cout => N_19293,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_1_RNITUGI4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_2_RNIJDE02: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNILU8P_14_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(14),
cin => N_19294);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_9_TRFWWBASICCELL_TEMP2_RNIV9EK8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD3\,
cout => N_19295,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_1_RNIF0M74: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_1_RNI778U1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNION6S_15_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(15),
cin => N_19296);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_10_TRFWWBASICCELL_TEMP2_RNINUSR8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD3\,
cout => N_19297,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_2_RNI06G74: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_RNIT2DM1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI915K_16_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(16),
cin => N_19298);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_11_TRFWWBASICCELL_TEMP2_RNI4J5P8: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD3\,
cout => N_19299,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_2_RNIVOU74: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_3_RNIML4R1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIT92I_17_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(17),
cin => N_19300);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_12_TRFWWBASICCELL_TEMP2_1_RNIF46C9: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD3\,
cout => N_19301,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_2_RNIC56C4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_1_RNIRUTJ1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIFFAL_18_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(18),
cin => N_19302);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_13_TRFWWBASICCELL_TEMP2_1_RNIN1F1A: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD3\,
cout => N_19303,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_3_RNIP7OH4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_1_RNI2BES1: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNI3STN_19_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(19),
cin => N_19304);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_14_TRFWWBASICCELL_TEMP2_RNIMEBFA: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD3\,
cout => N_19305,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD2\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(3),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_2\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_15_TRFWWBASICCELL_TEMP2_3_RNIJBHU4: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD2\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD1\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(2),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_1\);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_TRFWWRRAY_REMWTAGE57_16_TRFWWBASICCELL_TEMP2_1_RNI6AI62: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD1\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD0\,
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(1),
cin => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_0\);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_C_DPXX_CTRLXERSHFT_SUMIN_5_RNIL4TQ_20_\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "cin",
    lut_mask => "1001011011101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD0\,
cout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_CARRY_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_V\(0),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.CTRLXERSHFT.SUMIN_5\(20),
cin => N_19306);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_47\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_47\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000110010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100110101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111100110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_26\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011100010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_26\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_17\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_17\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000101010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100100100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100100001110110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100011001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100111111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_0_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_0_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_45\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_45\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000011101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101010101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_33\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101000101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_33\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111111010111110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011111010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_26\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_26\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110101011101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_20\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_20\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_11\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000010101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000111100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000111100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000010100101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010000010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_1_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_1_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111101110111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010111101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_49\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_49\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010011101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010111101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100111010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_33\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100101010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_33\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010111010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101110101011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001111000011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010110110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010110111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010011100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010011100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000101010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_2_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_2_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_61\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011101010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_61\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011111110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_47\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_47\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011101010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011111010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_38\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010001010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_38\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_37\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010101100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_37\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_33\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_33\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001010000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010010011010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010011011000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011001000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000110010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001110000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011111010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_3_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_3_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_61\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010100010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_61\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_58\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_58\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100010000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100111111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000000001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_46\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_46\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000101010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000111010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_35\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_35\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100011100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_33\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_33\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_21\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_21\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101011101010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001000010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001000000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010101000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001011101000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001011101010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_4_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001000010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_4_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_61\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_61\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_60\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100100001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_60\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_59\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_59\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_58\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_58\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100100011001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000011000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101001001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_54\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101110111011001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_49\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_49\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110010000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010110000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_37\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_37\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000010010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_35\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_35\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010111011001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_31\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_31\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111111011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001110010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011101011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_19\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_19\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_16\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_16\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000011001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000010011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100011000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000101001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000101011100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000101001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_5_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000110010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_5_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110101001101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_54\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111001001100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001110110011001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000010000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_37\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000001011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_37\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111100011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001100001001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_19\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110001001100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_19\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000011101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000101000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000111001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_6_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_6_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_61\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110101011101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_61\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_59\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_59\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100100010101101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111100001001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101110101111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_49\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_49\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010101010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011101010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_37\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010101010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_37\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100000101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000110100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010100111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011100011001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001001101101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011100101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010101101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001010101001111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001000111100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_7_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011101110111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_7_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010110001001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001111010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100001011001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_54\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001001011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_53\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000110000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_53\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_52\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_52\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001110010110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_46\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_46\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010110110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100110001111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_32\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_32\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_31\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_31\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110110000011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000010001011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101000001110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100100000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000001110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_19\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_19\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_17\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_17\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110000111001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010000110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000010101001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000010101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000011001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101110010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001010000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000110010010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_8_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101110010111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_8_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_61\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_61\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_58\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_58\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000101011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000000011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_54\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101100101111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_49\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000101000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_49\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100100000000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_46\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_46\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000001010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000001101011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_41\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_41\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_35\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_35\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_31\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_31\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111010101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001001100100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101100001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001101100101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_15\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_15\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100101100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1101100101000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000100000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_11\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100100101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100101101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000101101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1110000000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110000000101010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010000101000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100001101110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111000100100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1111100101101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_9_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_9_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_54\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000100101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000100100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_32\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_32\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_31\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_31\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100000110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000110110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010100110110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_17\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_17\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011011000010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010000000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100100001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_11\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000001100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110100000110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110111001100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011100000110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011001100101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000100101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011100000110001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110011000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111001110101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_10_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_10_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_54\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100001000001001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000001001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000101000101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011001101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000111000101100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101011100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_24\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_24\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000111001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100010010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_11\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000110100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010010110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000110111010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000110111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010001001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000100011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010101011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000010101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000110111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000100111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_11_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_11_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000000000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000001000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110000100110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_54\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001001000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_54\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101011000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010101011000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010000001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101011000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011010100111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_33\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_33\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001011000001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101000000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000011000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110010000100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_17\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_17\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101111010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011101010000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000100000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_11\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000100000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000100010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000000001000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011101110010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101111010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001101110010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001101110010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011101110010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_12_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001101110010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_12_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000010001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000010001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000001000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101110101000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111111001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_36\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_36\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001000011000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001010001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111010101000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000010101000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101010111010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011011101010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000010111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110001010010101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001010111101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001010010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111111101111111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_13_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001010010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_13_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_57\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100100001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_57\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_55\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_55\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1010101110100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_48\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001000000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_48\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_44\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000110000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_44\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_35\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000100100011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_35\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011100110111011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_31\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000001000001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_31\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110001100001010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000100010010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1011100000110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111101000101001")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1001100000110011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_24\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1100001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_24\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "1000001000000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110110101101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100110100100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_12\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000100010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_12\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_11\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000010000110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100010001110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011100110001011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110100000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001110000100101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010110001011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011010110100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010010110101011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010010110000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011110110101111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010010100000000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_14_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010010000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_14_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_56\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000110100000010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_56\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_50\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100110110000111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_50\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_45\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010001000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_45\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_43\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000010000000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_43\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_42\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100010010000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_42\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_34\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110110100011010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_34\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_30\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010100100111000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_30\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_29\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100100110000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_29\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_28\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000011000100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_28\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_27\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000000101001100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_27\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_25\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001100011010100")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_25\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_22\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0000100000001000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_22\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_18\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_18\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_14\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101011011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_14\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_13\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0110001101000101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_13\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_11\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_11\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_10\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0001000000010000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_10\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_9\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011000001011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_9\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_8\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011101010010")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_8\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_7\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111000001011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_7\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_6\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0011001001001101")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_6\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_5\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101011110")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_5\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_4\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101011000010111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_4\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_3\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100001100010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_3\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_2\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0101001000010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_2\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_1\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0111011101011111")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_1\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0__ROM_0\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0100011000010011")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0__ROM_0\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datad => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_PCTRL_NEW_19_15_0_62__ROM\: cycloneiii_lcell_comb generic map (
     sum_lutc_input => "datac",
    lut_mask => "0010000000100000")
port map (
combout => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_15_0_62__ROM\,
dataa => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
datab => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
datac => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85));
N_27907 <= not N_49;
N_27908 <= not \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RET_3: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2\(6),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.EXPADDERSHFT.EXPYBUS_2_RETI\(6),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_29_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(29),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(33),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_30_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(30),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(32),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RET_2: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES\,
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.LEFTSHIFTERBL.UN20_NOTSLRES_RETI\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_31_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(31),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(31),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_32_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(32),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_15\(30),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RET_1: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1\,
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP1_RETI\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_11_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(11),
d => N_19146,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_13_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(13),
d => N_19147,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RET_0: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD\,
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_RETI\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_RET: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2\,
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.FAX.UN13_NOTXZYFROMD_REP2_RETI\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_63_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(63),
d => \GRLFPC20.COMB.V.I.RES_1\(63),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_59_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(59),
d => \GRLFPC20.FPI.OP2_X\(62),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD7\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_58_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(58),
d => \GRLFPC20.FPI.OP2_X\(61),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD6\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_57_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(57),
d => \GRLFPC20.FPI.OP2_X\(60),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD5\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_56_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(56),
d => \GRLFPC20.FPI.OP2_X\(59),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD4\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_55_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(55),
d => \GRLFPC20.FPI.OP2_X\(58),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD3\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_54_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(54),
d => \GRLFPC20.FPI.OP2_X\(57),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD2\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_53_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(53),
d => \GRLFPC20.FPI.OP2_X\(56),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD1\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_52_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(52),
d => \GRLFPC20.FPI.OP2_X\(55),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD0\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_51_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(51),
d => \GRLFPC20.FPI.OP2_X\(54),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_50_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(50),
d => \GRLFPC20.FPI.OP2_X\(53),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_49_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(49),
d => \GRLFPC20.FPI.OP2_X\(52),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_48_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(48),
d => \GRLFPC20.FPI.OP2_X\(51),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_47_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(47),
d => \GRLFPC20.FPI.OP2_X\(50),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_46_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(46),
d => \GRLFPC20.FPI.OP2_X\(49),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_45_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(45),
d => \GRLFPC20.FPI.OP2_X\(48),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_44_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(44),
d => \GRLFPC20.FPI.OP2_X\(47),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_43_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(43),
d => \GRLFPC20.FPI.OP2_X\(46),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_42_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(42),
d => \GRLFPC20.FPI.OP2_X\(45),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_41_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(41),
d => \GRLFPC20.FPI.OP2_X\(44),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_40_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(40),
d => \GRLFPC20.FPI.OP2_X\(43),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_39_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(39),
d => \GRLFPC20.FPI.OP2_X\(42),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_38_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(38),
d => \GRLFPC20.FPI.OP2_X\(41),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_37_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(37),
d => \GRLFPC20.FPI.OP2_X\(40),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_36_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(36),
d => \GRLFPC20.FPI.OP2_X\(39),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_35_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(35),
d => \GRLFPC20.FPI.OP2_X\(38),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_34_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(34),
d => \GRLFPC20.FPI.OP2_X\(37),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_33_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(33),
d => \GRLFPC20.FPI.OP2_X\(36),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_32_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(32),
d => \GRLFPC20.FPI.OP2_X\(35),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_31_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(31),
d => \GRLFPC20.FPI.OP2_X\(34),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_30_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(30),
d => \GRLFPC20.FPI.OP2_X\(33),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_RES_29_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(29),
d => \GRLFPC20.FPI.OP2_X\(32),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\,
sload => \GRLFPC20.COMB.UN2_HOLDN_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_116_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(116),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_117_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(117),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(119),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_118_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(118),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(120),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_119_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(119),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(121),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_120_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(120),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(122),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_121_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(121),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(123),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_122_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(122),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(124),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_123_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(123),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(125),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_124_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(124),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(126),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_125_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(125),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(127),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_126_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(126),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(128),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_127_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(127),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(129),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_128_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(128),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(130),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_129_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(129),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(131),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_130_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(130),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(132),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_131_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(131),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(133),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_132_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(132),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(134),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_133_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(133),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(135),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_134_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(134),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(136),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_135_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(135),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(137),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_136_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(136),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(138),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_137_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(137),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(139),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_138_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(138),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(140),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_139_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(139),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_140_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(140),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_143_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(143),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(145),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_144_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(144),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(146),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_145_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(145),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(147),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_146_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(146),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(148),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_147_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(147),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(149),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_148_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(148),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(150),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_149_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(149),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(151),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_150_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(150),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(152),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_151_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(151),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(153),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_152_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(152),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(154),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_153_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(153),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(155),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_154_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(154),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(156),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_155_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(155),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(157),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_156_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(156),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(158),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_157_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(157),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(159),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_158_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(158),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(160),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_159_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(159),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(161),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_160_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(160),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(162),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_161_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(161),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(163),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_162_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(162),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(164),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_163_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(163),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(165),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_164_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(164),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(166),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_165_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(165),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(167),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_166_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(166),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(168),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_167_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(167),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(169),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_168_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(168),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(170),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_169_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(169),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_170_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(170),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.G_778\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_247_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(247),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(247),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_248_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(248),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(248),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_249_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(249),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(249),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_250_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(250),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(250),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_251_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(251),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(251),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_252_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(252),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(252),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_253_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(253),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(253),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_254_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(254),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(254),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_255_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(255),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(255),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_256_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(256),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(256),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_257_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(257),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(257),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.EXPBREGLOADEN\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_I_V: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.V\,
d => \GRLFPC20.R.I.V_1_0_G3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.V_1_0_G0_0\,
sclr => N_1_I,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_16_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(16),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_SCTRL_NEW_0_0__G0_I_M2\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_15_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(15),
d => N_27908,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_14_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(14),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_I_0_0__G0_0_M2\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_13_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(13),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_38_IV_I_0_0__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_12_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(12),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_R.SCTRL_39_IV\(0),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_11_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(11),
d => N_27907,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_10_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(10),
d => N_19148,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_9_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(9),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.UN17_U_RDN_I_0_503_I_A2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_8_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(8),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.U_RDN_1_520\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.RNDMODESELECT.TEMP\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_7_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(7),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_0_7__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_6_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(6),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(6),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(5),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.UN53_SCTRL_NEW\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(4),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(4),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(3),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW\(3),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(2),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_4_0_2__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(1),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_5_0_1__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_SCTRL_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.SCTRL\(0),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.SXC.SCTRL_NEW_6_0_0__G0_0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_85_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(85),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_0__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_84_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(84),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_1__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_83_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(83),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_2__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_82_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(82),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_0_3__G0_0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_81_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(81),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_4__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_80_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(80),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_5__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_79_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(79),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_6__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_78_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.MULTIPLEXORMULXFF.RESULT_1_IV_I_0_7__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_77_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(77),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW\(77),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_76_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(76),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN33_PCTRL_NEW_I_0_G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_74_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(74),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_18_0_74__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_73_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(73),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.STARTSHFT.UN3_NOTRESETORUNIMP\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_72_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(72),
d => N_19149,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_71_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(71),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.UN38_PCTRL_NEW_I_0_G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_70_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(70),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_69_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(69),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G2_0_529\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_11_0_69__G0_I_O4\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_68_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(68),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_65__G3\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_67_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(67),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_6_0_67__G3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_6_0_67__G0_E_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_66_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(66),
d => \GRLFPC20.FPI.START\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_65_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(65),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.PXS.PCTRL_NEW_2_0_65__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_64_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(64),
d => \GRLFPC20.FPI.RST_0_G0_X\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_63_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(63),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(0),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(0),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_62_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(62),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(1),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(1),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_61_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(61),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(2),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(2),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_60_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(60),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(3),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(3),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_59_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(59),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(4),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(4),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_58_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(58),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(5),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(5),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_57_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(57),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(6),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(6),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_56_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(56),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(7),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(7),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_55_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(55),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(8),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(8),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_54_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(54),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(9),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(9),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_53_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(53),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(10),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(10),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_52_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(52),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(11),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(11),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_51_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(51),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(12),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(12),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_50_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(50),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(13),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(13),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_49_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(49),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(14),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(14),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_48_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(48),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(15),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(15),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_47_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(47),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(16),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(16),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_46_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(46),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_46__G2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_45_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(45),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(18),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(18),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_44_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(44),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(19),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7_0_A2\(19),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_43_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(43),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(20),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(20),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_42_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(42),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(21),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(21),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_41_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(41),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_41__G4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_21_0_41__G3\,
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_40_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(40),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(23),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(23),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_39_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(39),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(24),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(24),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_38_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(38),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(25),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(25),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_36_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(36),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(26),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(26),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_35_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(35),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(27),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(27),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_34_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(34),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(28),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(28),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_33_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(33),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(29),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(29),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_28_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(28),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(34),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(34),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_27_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(27),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(35),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(35),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_26_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(26),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(36),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(36),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_25_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(25),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(37),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(37),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_24_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(24),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(38),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(38),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_23_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(23),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(39),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(39),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_22_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(22),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(40),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(40),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_21_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(21),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_21__G2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_20_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(20),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_20__G2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_19_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(19),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(43),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(43),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_18_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(18),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(44),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(44),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_17_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(17),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(45),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(45),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_16_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(16),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(46),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(46),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_15_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(15),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(47),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(47),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_14_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(14),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(48),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(48),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_12_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(12),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(50),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(50),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_9_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(9),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_9__G4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_9__G3\,
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_8_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(8),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(54),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(54),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_7_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(7),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(55),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(55),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_6_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(6),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(56),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(56),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(5),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(57),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(57),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(4),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(58),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(58),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(3),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(59),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(59),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(2),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_2_0_9__G4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(60),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(1),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(54),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(61),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_PCTRL_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(0),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_14\(62),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UPDATE_1\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.PCTRL_NEW_19_MUX_7\(62),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78),
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_377_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(377),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN1_GRFPUF_0\(0),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_376_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(376),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_DIVMULTV\(0),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_375_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(375),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_375__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_374_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(374),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_374__G0_0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_373_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(373),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN2_MIXOIN_25\(0),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_372_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(372),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(113),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_371_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(371),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(112),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_370_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(370),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(111),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_369_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(369),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(110),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_368_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(368),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(109),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_367_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(367),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(108),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_366_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(366),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(107),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_365_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(365),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(106),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_364_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(364),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(105),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_363_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(363),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(104),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_362_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(362),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(103),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_361_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(361),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(102),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_360_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(360),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(101),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_359_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(359),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(100),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_358_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(358),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(99),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_357_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(357),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(98),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_356_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(356),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(97),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_355_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(355),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(96),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_354_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(354),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(95),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_353_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(353),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(94),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_352_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(352),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(93),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_351_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(351),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(92),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_350_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(350),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(91),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_349_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(349),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(90),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_348_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(348),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(89),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_347_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(347),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(88),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_346_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(346),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(87),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_345_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(345),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(86),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_344_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(344),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(85),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_343_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(343),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(84),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_342_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(342),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(83),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_341_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(341),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(82),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_340_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(340),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(81),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_339_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(339),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(80),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_338_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(338),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(79),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_337_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(337),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(78),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_336_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(336),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(77),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_335_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(335),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(76),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_334_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(334),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(75),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_333_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(333),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(74),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_332_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(332),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(73),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_331_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(331),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(72),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_330_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(330),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(71),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_329_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(329),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(70),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_328_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(328),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(69),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_327_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(327),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(68),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_326_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(326),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(67),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_325_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(325),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(66),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_324_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(324),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(65),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_323_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(323),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(64),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_322_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(322),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(63),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_321_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(321),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(62),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_320_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(320),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23\(61),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_319_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(319),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_319__G3_0_X2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_318_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(318),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_318__G3_0_X2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_317_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(317),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.CO0\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_316_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(316),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_316__G3_0_X2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_315_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(315),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_315__G3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_314_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(314),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.3.CI_55_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_313_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(313),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.4.CI_54_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_312_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(312),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.5.CI_53_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_311_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(311),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.6.CI_52_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_310_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(310),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.7.CI_51_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_309_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(309),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.8.CI_50_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_308_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(308),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.9.CI_49_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_307_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(307),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.10.CI_48_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_306_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(306),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.11.CI_47_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_305_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(305),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.12.CI_46_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_304_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(304),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.13.CI_45_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_303_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(303),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.14.CI_44_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_302_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(302),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.15.CI_43_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_301_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(301),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.16.CI_42_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_300_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(300),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.17.CI_41_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_299_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(299),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.18.CI_40_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_298_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(298),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.19.CI_39_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_297_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(297),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.20.CI_38_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_296_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(296),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.21.CI_37_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_295_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(295),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.22.CI_36_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_294_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(294),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.23.CI_35_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_293_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(293),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.24.CI_34_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_292_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(292),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.25.CI_33_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_291_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(291),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.26.CI_32_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_290_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(290),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.27.CI_31_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_289_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(289),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.28.CI_30_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_288_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(288),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.29.CI_29_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_287_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(287),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.30.CI_28_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_286_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(286),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.31.CI_27_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_285_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(285),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.32.CI_26_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_284_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(284),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.33.CI_25_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_283_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(283),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.34.CI_24_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_282_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(282),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.35.CI_23_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_281_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(281),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.36.CI_22_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_280_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(280),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.37.CI_21_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_279_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(279),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.38.CI_20_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_278_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(278),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.39.CI_19_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_277_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(277),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.40.CI_18_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_276_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(276),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.41.CI_17_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_275_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(275),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.42.CI_16_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_274_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(274),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.43.CI_15_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_273_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(273),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.44.CI_14_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_272_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(272),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.45.CI_13_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_271_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(271),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.46.CI_12_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_270_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(270),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.47.CI_11_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_269_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(269),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.48.CI_10_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_268_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(268),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.49.CI_9_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_267_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(267),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.50.CI_8_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_266_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(266),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.51.CI_7_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_265_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(265),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.52.CI_6_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_264_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(264),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.53.CI_5_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_263_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(263),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.CI_4_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_262_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(262),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0\(0),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_261_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(261),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.TRFWWRRAY.54.SI_117_SUM1\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_260_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(260),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_23_1.SUM_0_A2\(0),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_259_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(259),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_8_1.SUM_0_A2\(0),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_258_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(258),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_258__G3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.UN2_NOTABORTWB\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_246_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(246),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(246),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_245_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(245),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(245),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_244_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(244),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(244),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_243_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(243),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(243),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_242_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(242),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(242),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_241_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(241),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(241),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_240_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(240),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(240),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_239_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(239),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(239),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_238_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(238),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(238),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_237_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(237),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(237),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_236_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(236),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(236),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_235_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(235),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(235),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_234_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(234),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(234),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_233_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(233),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(233),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_232_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(232),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(232),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_231_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(231),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD0\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_230_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(230),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD1\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_229_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(229),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_228_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(228),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_227_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(227),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_226_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(226),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_225_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(225),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_224_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(224),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_223_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(223),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_222_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(222),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_221_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(221),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_220_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(220),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_219_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(219),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_218_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(218),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_217_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(217),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_216_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(216),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_215_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(215),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_214_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(214),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_213_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(213),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_212_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(212),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_211_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(211),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_210_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(210),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_209_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(209),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_208_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(208),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_207_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(207),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_206_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(206),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_205_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(205),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_204_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(204),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_203_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(203),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_202_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(202),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_201_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(201),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_200_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(200),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_199_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(199),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD32\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_198_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(198),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD33\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_197_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(197),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD34\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_196_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(196),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD35\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_195_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(195),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD36\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_194_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(194),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD37\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_193_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(193),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD38\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_192_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(192),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD39\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_191_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(191),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD40\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_190_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(190),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD41\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_189_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(189),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD42\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_188_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(188),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD43\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_187_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(187),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD44\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_186_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(186),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD45\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_185_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(185),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD46\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_184_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(184),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD47\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_183_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(183),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD48\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_182_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(182),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD49\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_181_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(181),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD50\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_180_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(180),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD51\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_179_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(179),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD52\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_178_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(178),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD53\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_177_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(177),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD54\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_176_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(176),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD55\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_175_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(175),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD56\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_174_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(174),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD57\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_174__G2_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_173_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(173),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_173__G0_I\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_172_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(172),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_172__G0_0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_171_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(171),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(171),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_142_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(142),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(142),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_141_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(141),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(141),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_115_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(115),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(115),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_114_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(114),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_0_114__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_113_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(113),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(113),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_112_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(112),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_112__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_112__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_111_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(111),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_111__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_111__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_110_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(110),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_110__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_110__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_109_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(109),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_109__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_109__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_108_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(108),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_108__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_108__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_107_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(107),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_107__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_107__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_106_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(106),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_106__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_106__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_105_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(105),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_105__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_105__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_104_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(104),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_104__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_104__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_103_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(103),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_103__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_103__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_102_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(102),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_102__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_102__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_101_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(101),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_101__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_101__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_100_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(100),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_100__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_100__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_99_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(99),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_99__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_99__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_98_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(98),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_98__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_98__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_97_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(97),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_97__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_97__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_96_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(96),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_96__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_96__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_95_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(95),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_95__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_95__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_94_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(94),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_94__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_94__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_93_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(93),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_93__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_93__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_92_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(92),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_92__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_92__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_91_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(91),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_91__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_91__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_90_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(90),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_90__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_90__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_89_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(89),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_89__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_89__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_88_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(88),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_88__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_88__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_87_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(87),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_87__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_87__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_86_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(86),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_86__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_86__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_85_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(85),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_85__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_85__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_84_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(84),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_84__G2_X\,
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_0_84__G1\,
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_83_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(83),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_X\(83),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(83),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_82_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(82),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_X\(82),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(82),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_81_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(81),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19_X\(81),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(81),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_80_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(80),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(80),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(80),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_79_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(79),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(79),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(79),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_78_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(78),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(78),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(78),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_77_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(77),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(77),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(77),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_76_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(76),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(76),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(76),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_75_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(75),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(75),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(75),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_74_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(74),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(74),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(74),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_73_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(73),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(73),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(73),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_72_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(72),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(72),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(72),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_71_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(71),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(71),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(71),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_70_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(70),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(70),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(70),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_69_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(69),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(69),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(69),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_68_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(68),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(68),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(68),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_67_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(67),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(67),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(67),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_66_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(66),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(66),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(66),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_65_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(65),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(65),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(65),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_64_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(64),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(64),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(64),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_63_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(63),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(63),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(63),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_62_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(62),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(62),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(62),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_61_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(61),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.DPATH_NEW_19\(61),
clk => N_2,
clrn => VCC,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_M3\(61),
sload => \GRLFPC20.FPI.LDOP_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_60_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(60),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(60),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_59_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(59),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(59),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_58_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(58),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH\(58),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_57_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(57),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(57),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(57),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_56_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(56),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(56),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(56),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_55_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(55),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(55),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(55),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_54_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(54),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(54),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(54),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_53_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(53),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(53),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(53),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_52_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(52),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(52),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(52),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_51_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(51),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(51),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(51),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_50_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(50),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(50),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(50),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_49_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(49),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(49),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(49),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_48_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(48),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(48),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(48),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_47_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(47),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(47),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(47),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_46_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(46),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(46),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(46),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_45_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(45),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(45),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(45),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_44_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(44),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(44),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(44),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_43_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(43),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(43),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(43),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_42_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(42),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(42),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(42),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_41_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(41),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(41),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(41),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_40_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(40),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(40),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(40),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_39_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(39),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(39),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(39),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_38_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(38),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(38),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(38),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_37_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(37),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(37),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(37),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_36_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(36),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(36),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(36),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_35_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(35),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(35),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(35),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_34_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(34),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(34),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(34),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_33_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(33),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(33),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(33),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_32_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(32),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(32),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(32),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_31_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(31),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(31),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(31),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_30_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(30),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(30),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(30),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_29_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(29),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(29),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(29),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_28_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(28),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(28),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(28),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_27_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(27),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(27),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(27),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_26_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(26),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(26),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(26),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_25_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(25),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(25),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(25),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_24_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(24),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(24),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(24),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_23_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(23),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(23),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(23),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_22_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(22),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(22),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(22),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_21_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(21),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(21),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(21),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_20_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(20),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(20),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(20),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_19_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(19),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(19),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(19),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_18_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(18),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(18),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(18),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_17_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(17),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(17),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(17),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_16_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(16),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(16),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(16),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_15_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(15),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(15),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(15),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_14_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(14),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(14),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(14),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_13_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(13),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(13),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(13),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_12_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(12),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(12),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(12),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_11_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(11),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(11),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(11),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_10_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(10),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(10),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(10),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_9_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(9),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(9),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(9),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_8_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(8),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(8),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(8),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_7_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(7),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(7),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(7),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_6_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(6),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(6),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(6),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(5),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(5),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(5),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(4),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(4),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(4),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(3),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(3),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(3),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(2),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(2),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(2),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(1),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(1),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(1),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_GRFPUL_GEN0_GRLFPU0_R_DPATH_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.DPATH\(0),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_4\(0),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.C.DPXX.XZAREGLOADEN\,
asdata => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_5\(0),
sload => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
GRLFPC20_R_MK_HOLDN2: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.MK.HOLDN2\,
d => \GRLFPC20.R.MK.HOLDN1\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_MK_RST: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.MK.RST\,
d => \GRLFPC20.COMB.V.MK.RST_1_0_G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_MK_RST2: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.MK.RST2\,
d => \GRLFPC20.R.MK.RST\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_MK_LDOP: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.MK.LDOP\,
d => \GRLFPC20.RIN.MK.LDOP_X\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_X_RDD_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.X.RDD\(0),
d => \GRLFPC20.R.M.RDD\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_M_RDD_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.M.RDD\(0),
d => \GRLFPC20.R.E.RDD\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_E_RDD_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.E.RDD\(0),
d => \GRLFPC20.R.A.RDD\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RDD_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RDD\(0),
d => \GRLFPC20.R.A.RDD_0_0_0__G1_0\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_X_SEQERR_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.X.SEQERR\(0),
d => \GRLFPC20.R.M.SEQERR\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_M_SEQERR_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.M.SEQERR\(0),
d => \GRLFPC20.R.E.SEQERR\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_E_SEQERR_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.E.SEQERR\(0),
d => \GRLFPC20.R.A.SEQERR\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_SEQERR_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.SEQERR\(0),
d => \GRLFPC20.R.A.SEQERR_0_0_0__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_I_EXEC: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.EXEC\,
d => \GRLFPC20.R.I.EXEC_0_0_G1_0_549_I\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_ST: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.ST\,
d => \GRLFPC20.R.A.ST_0_0_G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_LD: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.LD\,
d => \GRLFPC20.R.A.LD_0_0_G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_FPOP: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.FPOP\,
d => \GRLFPC20.R.A.FPOP_0_0_G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_AFSR: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.AFSR\,
d => \GRLFPC20.R.A.AFSR_0_0_G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_AFQ: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.AFQ\,
d => \GRLFPC20.R.A.AFQ_0_0_G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_RS1D: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS1D\,
d => \GRLFPC20.COMB.RS1D_1_U\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_RS2D: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS2D\,
d => \GRLFPC20.COMB.RS2D_1_IV\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_FSR_NONSTD: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.NONSTD\,
d => \GRLFPC20.R.FSR.NONSTD_0_0_G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_418,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
GRLFPC20_R_I_RDD: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RDD\,
d => \GRLFPC20.R.I.RDD_0_0_G1_0_574_I\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_A_MOV: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.MOV\,
d => \GRLFPC20.R.A.MOV_0_0_G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_X_LD: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.X.LD\,
d => \GRLFPC20.R.X.LD_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_X_FPOP: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.X.FPOP\,
d => \GRLFPC20.R.X.FPOP_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_X_AFSR: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.X.AFSR\,
d => \GRLFPC20.R.X.AFSR_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_X_AFQ: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.X.AFQ\,
d => \GRLFPC20.R.X.AFQ_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_M_LD: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.M.LD\,
d => \GRLFPC20.R.M.LD_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_M_FPOP: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.M.FPOP\,
d => \GRLFPC20.R.M.FPOP_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_M_AFSR: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.M.AFSR\,
d => \GRLFPC20.R.M.AFSR_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_M_AFQ: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.M.AFQ\,
d => \GRLFPC20.R.M.AFQ_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_E_LD: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.E.LD\,
d => \GRLFPC20.R.E.LD_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_E_FPOP: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.E.FPOP\,
d => \GRLFPC20.R.E.FPOP_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_E_AFSR: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.E.AFSR\,
d => \GRLFPC20.R.E.AFSR_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_E_AFQ: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.E.AFQ\,
d => \GRLFPC20.R.E.AFQ_0_0_G1_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_MK_HOLDN1: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.MK.HOLDN1\,
d => \GRLFPC20.R.MK.HOLDN1_0_0_G0_X\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_MK_BUSY: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.MK.BUSY\,
d => \GRLFPC20.R.MK.BUSY_0_0_G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
GRLFPC20_R_MK_BUSY2: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.MK.BUSY2\,
d => \GRLFPC20.R.MK.BUSY2_0_0_G0_X\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(2),
d => N_289,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(3),
d => N_290,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(4),
d => N_291,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(5),
d => N_292,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_6_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(6),
d => N_293,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_7_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(7),
d => N_294,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_8_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(8),
d => N_295,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_9_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(9),
d => N_296,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_10_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(10),
d => N_297,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_11_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(11),
d => N_298,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_12_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(12),
d => N_299,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_13_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(13),
d => N_300,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_14_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(14),
d => N_301,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_15_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(15),
d => N_302,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_16_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(16),
d => N_303,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_17_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(17),
d => N_304,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_18_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(18),
d => N_305,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_19_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(19),
d => N_306,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_20_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(20),
d => N_307,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_21_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(21),
d => N_308,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_22_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(22),
d => N_309,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_23_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(23),
d => N_310,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_24_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(24),
d => N_311,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_25_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(25),
d => N_312,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_26_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(26),
d => N_313,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_27_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(27),
d => N_314,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_28_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(28),
d => N_315,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_29_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(29),
d => N_316,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_30_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(30),
d => N_317,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_PC_31_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.PC\(31),
d => N_318,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.I.PC_1_0_2__G2_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_CC_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.CC\(0),
d => \GRLFPC20.R.I.CC_0_0_0__G4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_CC_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.CC\(1),
d => \GRLFPC20.R.I.CC_0_0_1__G4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_E_STDATA_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(0),
d => \GRLFPC20.R.E.STDATA_1_0_0__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_0__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(1),
d => \GRLFPC20.R.E.STDATA_1_0_1__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_1__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(2),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(2),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(2),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(3),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(3),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(3),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(4),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(4),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(4),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(5),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(5),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(5),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_6_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(6),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(6),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(6),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_7_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(7),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(7),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(7),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_8_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(8),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(8),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(8),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_9_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(9),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(9),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(9),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_10_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(10),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(10),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(10),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_11_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(11),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(11),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(11),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_12_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(12),
d => \GRLFPC20.R.E.STDATA_1_0_12__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_12__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_13_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(13),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(13),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(13),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_14_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(14),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(14),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(14),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_15_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(15),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(15),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(15),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_16_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(16),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(16),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(16),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_17_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(17),
d => \GRLFPC20.R.E.STDATA_1_0_17__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_17__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_18_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(18),
d => \GRLFPC20.R.E.STDATA_1_0_18__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_18__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_19_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(19),
d => \GRLFPC20.R.E.STDATA_1_0_19__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_19__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_20_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(20),
d => \GRLFPC20.R.E.STDATA_1_0_20__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_20__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_21_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(21),
d => \GRLFPC20.R.E.STDATA_1_0_21__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_21__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_22_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(22),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(22),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(22),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_23_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(23),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(23),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(23),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_24_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(24),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(24),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(24),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_25_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(25),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(25),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(25),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_26_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(26),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(26),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(26),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_27_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(27),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(27),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(27),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_28_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(28),
d => \GRLFPC20.R.E.STDATA_1_0_28__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_28__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_29_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(29),
d => \GRLFPC20.R.E.STDATA_1_0_29__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.E.STDATA_1_0_29__G2\,
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_30_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(30),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(30),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(30),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_E_STDATA_31_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_DATAZ(31),
d => \GRLFPC20.COMB.V.E.STDATA_1_0_X\(31),
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.COMB.V.E.STDATA_1_1\(31),
sload => \GRLFPC20.R.A.AFQ_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND,
	sclr => GND);
\GRLFPC20_R_I_INST_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(0),
d => N_319,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(0),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(1),
d => N_320,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(1),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(2),
d => N_321,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(2),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(3),
d => N_322,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(3),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(4),
d => N_323,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(4),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(5),
d => N_324,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(5),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_6_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(6),
d => N_325,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(6),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_7_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(7),
d => N_326,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(7),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_8_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(8),
d => N_327,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(8),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_9_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(9),
d => N_328,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(9),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_10_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(10),
d => N_329,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(10),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_11_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(11),
d => N_330,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(11),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_12_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(12),
d => N_331,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(12),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_13_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(13),
d => N_332,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(13),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_14_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(14),
d => N_333,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(14),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_15_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(15),
d => N_334,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(15),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_16_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(16),
d => N_335,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(16),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_17_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(17),
d => N_336,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(17),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_18_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(18),
d => N_337,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(18),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_19_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(19),
d => N_338,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(19),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_20_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(20),
d => N_339,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(20),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_21_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(21),
d => N_340,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(21),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_22_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(22),
d => N_341,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(22),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_23_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(23),
d => N_342,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(23),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_24_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(24),
d => N_343,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(24),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_25_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(25),
d => N_344,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(25),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_26_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(26),
d => N_345,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(26),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_27_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(27),
d => N_346,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(27),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_28_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(28),
d => N_347,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(28),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_29_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(29),
d => N_348,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(29),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_30_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(30),
d => N_349,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(30),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_I_INST_31_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.INST\(31),
d => N_350,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => \GRLFPC20.R.I.INST\(31),
sclr => N_1_I,
sload => \GRLFPC20.V.I.EXEC_0_SQMUXA_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_FSR_RD_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.RD\(0),
d => \GRLFPC20.R.FSR.RD_0_0_0__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_426,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_FSR_RD_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.RD\(1),
d => \GRLFPC20.R.FSR.RD_0_0_1__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_427,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_FSR_TEM_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.TEM\(0),
d => \GRLFPC20.R.FSR.TEM_1_0_0__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_419,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_FSR_TEM_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.TEM\(1),
d => \GRLFPC20.R.FSR.TEM_1_0_1__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_420,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_FSR_TEM_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.TEM\(2),
d => \GRLFPC20.R.FSR.TEM_1_0_2__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_421,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_FSR_TEM_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.TEM\(3),
d => \GRLFPC20.R.FSR.TEM_1_0_3__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_422,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_FSR_TEM_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.TEM\(4),
d => \GRLFPC20.R.FSR.TEM_1_0_4__G3_X\,
clk => N_2,
clrn => VCC,
ena => N_3,
asdata => N_423,
sclr => N_1_I,
sload => \GRLFPC20.V.STATE_0_SQMUXA_1_X_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	aload => GND);
\GRLFPC20_R_STATE_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.STATE\(0),
d => \GRLFPC20.R.STATE_0_0_0__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_STATE_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.STATE\(1),
d => \GRLFPC20.R.STATE_0_0_1__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_FTT_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.FTT\(0),
d => \GRLFPC20.R.FSR.FTT_1_0_0__G2_0_600_I\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.FSR.FTT_1_0_0__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_FTT_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.FTT\(1),
d => \GRLFPC20.R.FSR.FTT_1_0_1__G2_0_624_I\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.FSR.FTT_1_0_0__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_FTT_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.FTT\(2),
d => \GRLFPC20.R.FSR.FTT_1_0_2__G2\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.R.FSR.FTT_1_0_0__G0_I_O4_I\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RF1REN_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RF1REN\(2),
d => \GRLFPC20.COMB.V.A.RF1REN_1\(2),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RF1REN_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RF1REN\(1),
d => \GRLFPC20.COMB.V.A.RF1REN_1_670_I\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RF2REN_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RF2REN\(2),
d => \GRLFPC20.COMB.V.A.RF2REN_1_0_701_I\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RF2REN_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RF2REN\(1),
d => \GRLFPC20.COMB.V.A.RF2REN_1_734_I\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_FCC_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_CCZ(0),
d => \GRLFPC20.COMB.V.FSR.FCC_1\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_FCC_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => CPO_CCZ(1),
d => \GRLFPC20.COMB.V.FSR.FCC_1\(1),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_AEXC_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.AEXC\(0),
d => \GRLFPC20.R.FSR.AEXC_1_0_0__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_AEXC_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.AEXC\(1),
d => \GRLFPC20.R.FSR.AEXC_1_0_1__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_AEXC_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.AEXC\(2),
d => \GRLFPC20.R.FSR.AEXC_1_0_2__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_AEXC_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.AEXC\(3),
d => \GRLFPC20.R.FSR.AEXC_1_0_3__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_AEXC_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.AEXC\(4),
d => \GRLFPC20.R.FSR.AEXC_1_0_4__G1\,
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_CEXC_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.CEXC\(0),
d => \GRLFPC20.COMB.V.FSR.CEXC_1\(0),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_CEXC_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.CEXC\(1),
d => \GRLFPC20.COMB.V.FSR.CEXC_1\(1),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_CEXC_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.CEXC\(2),
d => \GRLFPC20.COMB.V.FSR.CEXC_1\(2),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_CEXC_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.CEXC\(3),
d => \GRLFPC20.COMB.V.FSR.CEXC_1\(3),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_FSR_CEXC_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.FSR.CEXC\(4),
d => \GRLFPC20.COMB.V.FSR.CEXC_1\(4),
clk => N_2,
clrn => VCC,
ena => N_3,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_EXC_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.EXC\(0),
d => \GRLFPC20.R.I.EXC_2_0_0__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_EXC_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.EXC\(1),
d => \GRLFPC20.R.I.EXC_0\(1),
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_EXC_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.EXC\(2),
d => \GRLFPC20.R.I.EXC_2_0_2__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_EXC_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.EXC\(3),
d => \GRLFPC20.R.I.EXC_2_0_3__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_EXC_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.EXC\(4),
d => \GRLFPC20.R.I.EXC_2_0_4__G3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.G_884\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_EXC_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.EXC\(5),
d => \GRLFPC20.R.I.EXC_2_0_5__G0\,
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS1_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS1\(0),
d => \GRLFPC20.COMB.RS1_1\(0),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS1_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS1\(1),
d => \GRLFPC20.COMB.RS1_1\(1),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS1_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS1\(2),
d => \GRLFPC20.COMB.RS1_1\(2),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS1_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS1\(3),
d => \GRLFPC20.COMB.RS1_1\(3),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS1_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS1\(4),
d => \GRLFPC20.COMB.RS1_1\(4),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(0),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD3\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(1),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD4\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(2),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD5\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(3),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD6\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(4),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD7\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_5_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(5),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD8\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_6_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(6),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD9\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_7_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(7),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD10\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_8_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(8),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD11\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_9_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(9),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD12\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_10_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(10),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD13\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_11_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(11),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD14\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_12_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(12),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD15\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_13_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(13),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD16\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_14_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(14),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD17\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_15_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(15),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD18\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_16_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(16),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD19\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_17_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(17),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD20\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_18_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(18),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD21\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_19_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(19),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD22\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_20_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(20),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD23\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_21_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(21),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD24\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_22_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(22),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD25\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_23_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(23),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD26\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_24_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(24),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD27\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_25_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(25),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD28\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_26_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(26),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD29\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_27_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(27),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD30\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_28_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(28),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUF_ADD31\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_60_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(60),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD8\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_61_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(61),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD9\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_I_RES_62_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.I.RES\(62),
d => \GRLFPC20.GRFPUL_GEN0.GRLFPU0.UN6_GRFPUE_ADD10\,
clk => N_2,
clrn => VCC,
ena => \GRLFPC20.COMB.UN19_IUEXEC\,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS2_0_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS2\(0),
d => \GRLFPC20.COMB.RS2_1\(0),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS2_1_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS2\(1),
d => \GRLFPC20.COMB.RS2_1\(1),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS2_2_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS2\(2),
d => \GRLFPC20.COMB.RS2_1\(2),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS2_3_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS2\(3),
d => \GRLFPC20.COMB.RS2_1\(3),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
\GRLFPC20_R_A_RS2_4_\: dffeas generic map (
    is_wysiwyg => "true" )
port map (
q => \GRLFPC20.R.A.RS2\(4),
d => \GRLFPC20.COMB.RS2_1\(4),
clk => N_2,
clrn => VCC,
	devpor => devpor,
	devclrn => devclrn,
	prn => VCC,
	ena => VCC,
	asdata => GND,
	aload => GND,
	sclr => GND,
	sload => GND);
N_1 <= RST_INTERNAL;
N_2 <= CLK_INTERNAL;
N_3 <= HOLDN_INTERNAL;
N_4 <= CPI_FLUSH_INTERNAL;
N_5 <= CPI_EXACK_INTERNAL;
N_6 <= CPI_A_RS1_INTERNAL;
N_7 <= CPI_A_RS1_INTERNAL_0;
N_8 <= CPI_A_RS1_INTERNAL_1;
N_9 <= CPI_A_RS1_INTERNAL_2;
N_10 <= CPI_A_RS1_INTERNAL_3;
N_11 <= CPI_D_PC_INTERNAL;
N_12 <= CPI_D_PC_INTERNAL_0;
N_13 <= CPI_D_PC_INTERNAL_1;
N_14 <= CPI_D_PC_INTERNAL_2;
N_15 <= CPI_D_PC_INTERNAL_3;
N_16 <= CPI_D_PC_INTERNAL_4;
N_17 <= CPI_D_PC_INTERNAL_5;
N_18 <= CPI_D_PC_INTERNAL_6;
N_19 <= CPI_D_PC_INTERNAL_7;
N_20 <= CPI_D_PC_INTERNAL_8;
N_21 <= CPI_D_PC_INTERNAL_9;
N_22 <= CPI_D_PC_INTERNAL_10;
N_23 <= CPI_D_PC_INTERNAL_11;
N_24 <= CPI_D_PC_INTERNAL_12;
N_25 <= CPI_D_PC_INTERNAL_13;
N_26 <= CPI_D_PC_INTERNAL_14;
N_27 <= CPI_D_PC_INTERNAL_15;
N_28 <= CPI_D_PC_INTERNAL_16;
N_29 <= CPI_D_PC_INTERNAL_17;
N_30 <= CPI_D_PC_INTERNAL_18;
N_31 <= CPI_D_PC_INTERNAL_19;
N_32 <= CPI_D_PC_INTERNAL_20;
N_33 <= CPI_D_PC_INTERNAL_21;
N_34 <= CPI_D_PC_INTERNAL_22;
N_35 <= CPI_D_PC_INTERNAL_23;
N_36 <= CPI_D_PC_INTERNAL_24;
N_37 <= CPI_D_PC_INTERNAL_25;
N_38 <= CPI_D_PC_INTERNAL_26;
N_39 <= CPI_D_PC_INTERNAL_27;
N_40 <= CPI_D_PC_INTERNAL_28;
N_41 <= CPI_D_PC_INTERNAL_29;
N_42 <= CPI_D_PC_INTERNAL_30;
N_43 <= CPI_D_INST_INTERNAL;
N_44 <= CPI_D_INST_INTERNAL_0;
N_45 <= CPI_D_INST_INTERNAL_1;
N_46 <= CPI_D_INST_INTERNAL_2;
N_47 <= CPI_D_INST_INTERNAL_3;
N_48 <= CPI_D_INST_INTERNAL_4;
N_49 <= CPI_D_INST_INTERNAL_5;
N_50 <= CPI_D_INST_INTERNAL_6;
N_51 <= CPI_D_INST_INTERNAL_7;
N_52 <= CPI_D_INST_INTERNAL_8;
N_53 <= CPI_D_INST_INTERNAL_9;
N_54 <= CPI_D_INST_INTERNAL_10;
N_55 <= CPI_D_INST_INTERNAL_11;
N_56 <= CPI_D_INST_INTERNAL_12;
N_57 <= CPI_D_INST_INTERNAL_13;
N_58 <= CPI_D_INST_INTERNAL_14;
N_59 <= CPI_D_INST_INTERNAL_15;
N_60 <= CPI_D_INST_INTERNAL_16;
N_61 <= CPI_D_INST_INTERNAL_17;
N_62 <= CPI_D_INST_INTERNAL_18;
N_63 <= CPI_D_INST_INTERNAL_19;
N_64 <= CPI_D_INST_INTERNAL_20;
N_65 <= CPI_D_INST_INTERNAL_21;
N_66 <= CPI_D_INST_INTERNAL_22;
N_67 <= CPI_D_INST_INTERNAL_23;
N_68 <= CPI_D_INST_INTERNAL_24;
N_69 <= CPI_D_INST_INTERNAL_25;
N_70 <= CPI_D_INST_INTERNAL_26;
N_71 <= CPI_D_INST_INTERNAL_27;
N_72 <= CPI_D_INST_INTERNAL_28;
N_73 <= CPI_D_INST_INTERNAL_29;
N_74 <= CPI_D_INST_INTERNAL_30;
N_75 <= CPI_D_CNT_INTERNAL;
N_76 <= CPI_D_CNT_INTERNAL_0;
N_77 <= CPI_D_TRAP_INTERNAL;
N_78 <= CPI_D_ANNUL_INTERNAL;
N_79 <= CPI_D_PV_INTERNAL;
N_80 <= CPI_A_PC_INTERNAL;
N_81 <= CPI_A_PC_INTERNAL_0;
N_82 <= CPI_A_PC_INTERNAL_1;
N_83 <= CPI_A_PC_INTERNAL_2;
N_84 <= CPI_A_PC_INTERNAL_3;
N_85 <= CPI_A_PC_INTERNAL_4;
N_86 <= CPI_A_PC_INTERNAL_5;
N_87 <= CPI_A_PC_INTERNAL_6;
N_88 <= CPI_A_PC_INTERNAL_7;
N_89 <= CPI_A_PC_INTERNAL_8;
N_90 <= CPI_A_PC_INTERNAL_9;
N_91 <= CPI_A_PC_INTERNAL_10;
N_92 <= CPI_A_PC_INTERNAL_11;
N_93 <= CPI_A_PC_INTERNAL_12;
N_94 <= CPI_A_PC_INTERNAL_13;
N_95 <= CPI_A_PC_INTERNAL_14;
N_96 <= CPI_A_PC_INTERNAL_15;
N_97 <= CPI_A_PC_INTERNAL_16;
N_98 <= CPI_A_PC_INTERNAL_17;
N_99 <= CPI_A_PC_INTERNAL_18;
N_100 <= CPI_A_PC_INTERNAL_19;
N_101 <= CPI_A_PC_INTERNAL_20;
N_102 <= CPI_A_PC_INTERNAL_21;
N_103 <= CPI_A_PC_INTERNAL_22;
N_104 <= CPI_A_PC_INTERNAL_23;
N_105 <= CPI_A_PC_INTERNAL_24;
N_106 <= CPI_A_PC_INTERNAL_25;
N_107 <= CPI_A_PC_INTERNAL_26;
N_108 <= CPI_A_PC_INTERNAL_27;
N_109 <= CPI_A_PC_INTERNAL_28;
N_110 <= CPI_A_PC_INTERNAL_29;
N_111 <= CPI_A_PC_INTERNAL_30;
N_112 <= CPI_A_INST_INTERNAL;
N_113 <= CPI_A_INST_INTERNAL_0;
N_114 <= CPI_A_INST_INTERNAL_1;
N_115 <= CPI_A_INST_INTERNAL_2;
N_116 <= CPI_A_INST_INTERNAL_3;
N_117 <= CPI_A_INST_INTERNAL_4;
N_118 <= CPI_A_INST_INTERNAL_5;
N_119 <= CPI_A_INST_INTERNAL_6;
N_120 <= CPI_A_INST_INTERNAL_7;
N_121 <= CPI_A_INST_INTERNAL_8;
N_122 <= CPI_A_INST_INTERNAL_9;
N_123 <= CPI_A_INST_INTERNAL_10;
N_124 <= CPI_A_INST_INTERNAL_11;
N_125 <= CPI_A_INST_INTERNAL_12;
N_126 <= CPI_A_INST_INTERNAL_13;
N_127 <= CPI_A_INST_INTERNAL_14;
N_128 <= CPI_A_INST_INTERNAL_15;
N_129 <= CPI_A_INST_INTERNAL_16;
N_130 <= CPI_A_INST_INTERNAL_17;
N_131 <= CPI_A_INST_INTERNAL_18;
N_132 <= CPI_A_INST_INTERNAL_19;
N_133 <= CPI_A_INST_INTERNAL_20;
N_134 <= CPI_A_INST_INTERNAL_21;
N_135 <= CPI_A_INST_INTERNAL_22;
N_136 <= CPI_A_INST_INTERNAL_23;
N_137 <= CPI_A_INST_INTERNAL_24;
N_138 <= CPI_A_INST_INTERNAL_25;
N_139 <= CPI_A_INST_INTERNAL_26;
N_140 <= CPI_A_INST_INTERNAL_27;
N_141 <= CPI_A_INST_INTERNAL_28;
N_142 <= CPI_A_INST_INTERNAL_29;
N_143 <= CPI_A_INST_INTERNAL_30;
N_144 <= CPI_A_CNT_INTERNAL;
N_145 <= CPI_A_CNT_INTERNAL_0;
N_146 <= CPI_A_TRAP_INTERNAL;
N_147 <= CPI_A_ANNUL_INTERNAL;
N_148 <= CPI_A_PV_INTERNAL;
N_149 <= CPI_E_PC_INTERNAL;
N_150 <= CPI_E_PC_INTERNAL_0;
N_151 <= CPI_E_PC_INTERNAL_1;
N_152 <= CPI_E_PC_INTERNAL_2;
N_153 <= CPI_E_PC_INTERNAL_3;
N_154 <= CPI_E_PC_INTERNAL_4;
N_155 <= CPI_E_PC_INTERNAL_5;
N_156 <= CPI_E_PC_INTERNAL_6;
N_157 <= CPI_E_PC_INTERNAL_7;
N_158 <= CPI_E_PC_INTERNAL_8;
N_159 <= CPI_E_PC_INTERNAL_9;
N_160 <= CPI_E_PC_INTERNAL_10;
N_161 <= CPI_E_PC_INTERNAL_11;
N_162 <= CPI_E_PC_INTERNAL_12;
N_163 <= CPI_E_PC_INTERNAL_13;
N_164 <= CPI_E_PC_INTERNAL_14;
N_165 <= CPI_E_PC_INTERNAL_15;
N_166 <= CPI_E_PC_INTERNAL_16;
N_167 <= CPI_E_PC_INTERNAL_17;
N_168 <= CPI_E_PC_INTERNAL_18;
N_169 <= CPI_E_PC_INTERNAL_19;
N_170 <= CPI_E_PC_INTERNAL_20;
N_171 <= CPI_E_PC_INTERNAL_21;
N_172 <= CPI_E_PC_INTERNAL_22;
N_173 <= CPI_E_PC_INTERNAL_23;
N_174 <= CPI_E_PC_INTERNAL_24;
N_175 <= CPI_E_PC_INTERNAL_25;
N_176 <= CPI_E_PC_INTERNAL_26;
N_177 <= CPI_E_PC_INTERNAL_27;
N_178 <= CPI_E_PC_INTERNAL_28;
N_179 <= CPI_E_PC_INTERNAL_29;
N_180 <= CPI_E_PC_INTERNAL_30;
N_181 <= CPI_E_INST_INTERNAL;
N_182 <= CPI_E_INST_INTERNAL_0;
N_183 <= CPI_E_INST_INTERNAL_1;
N_184 <= CPI_E_INST_INTERNAL_2;
N_185 <= CPI_E_INST_INTERNAL_3;
N_186 <= CPI_E_INST_INTERNAL_4;
N_187 <= CPI_E_INST_INTERNAL_5;
N_188 <= CPI_E_INST_INTERNAL_6;
N_189 <= CPI_E_INST_INTERNAL_7;
N_190 <= CPI_E_INST_INTERNAL_8;
N_191 <= CPI_E_INST_INTERNAL_9;
N_192 <= CPI_E_INST_INTERNAL_10;
N_193 <= CPI_E_INST_INTERNAL_11;
N_194 <= CPI_E_INST_INTERNAL_12;
N_195 <= CPI_E_INST_INTERNAL_13;
N_196 <= CPI_E_INST_INTERNAL_14;
N_197 <= CPI_E_INST_INTERNAL_15;
N_198 <= CPI_E_INST_INTERNAL_16;
N_199 <= CPI_E_INST_INTERNAL_17;
N_200 <= CPI_E_INST_INTERNAL_18;
N_201 <= CPI_E_INST_INTERNAL_19;
N_202 <= CPI_E_INST_INTERNAL_20;
N_203 <= CPI_E_INST_INTERNAL_21;
N_204 <= CPI_E_INST_INTERNAL_22;
N_205 <= CPI_E_INST_INTERNAL_23;
N_206 <= CPI_E_INST_INTERNAL_24;
N_207 <= CPI_E_INST_INTERNAL_25;
N_208 <= CPI_E_INST_INTERNAL_26;
N_209 <= CPI_E_INST_INTERNAL_27;
N_210 <= CPI_E_INST_INTERNAL_28;
N_211 <= CPI_E_INST_INTERNAL_29;
N_212 <= CPI_E_INST_INTERNAL_30;
N_213 <= CPI_E_CNT_INTERNAL;
N_214 <= CPI_E_CNT_INTERNAL_0;
N_215 <= CPI_E_TRAP_INTERNAL;
N_216 <= CPI_E_ANNUL_INTERNAL;
N_217 <= CPI_E_PV_INTERNAL;
N_218 <= CPI_M_PC_INTERNAL;
N_219 <= CPI_M_PC_INTERNAL_0;
N_220 <= CPI_M_PC_INTERNAL_1;
N_221 <= CPI_M_PC_INTERNAL_2;
N_222 <= CPI_M_PC_INTERNAL_3;
N_223 <= CPI_M_PC_INTERNAL_4;
N_224 <= CPI_M_PC_INTERNAL_5;
N_225 <= CPI_M_PC_INTERNAL_6;
N_226 <= CPI_M_PC_INTERNAL_7;
N_227 <= CPI_M_PC_INTERNAL_8;
N_228 <= CPI_M_PC_INTERNAL_9;
N_229 <= CPI_M_PC_INTERNAL_10;
N_230 <= CPI_M_PC_INTERNAL_11;
N_231 <= CPI_M_PC_INTERNAL_12;
N_232 <= CPI_M_PC_INTERNAL_13;
N_233 <= CPI_M_PC_INTERNAL_14;
N_234 <= CPI_M_PC_INTERNAL_15;
N_235 <= CPI_M_PC_INTERNAL_16;
N_236 <= CPI_M_PC_INTERNAL_17;
N_237 <= CPI_M_PC_INTERNAL_18;
N_238 <= CPI_M_PC_INTERNAL_19;
N_239 <= CPI_M_PC_INTERNAL_20;
N_240 <= CPI_M_PC_INTERNAL_21;
N_241 <= CPI_M_PC_INTERNAL_22;
N_242 <= CPI_M_PC_INTERNAL_23;
N_243 <= CPI_M_PC_INTERNAL_24;
N_244 <= CPI_M_PC_INTERNAL_25;
N_245 <= CPI_M_PC_INTERNAL_26;
N_246 <= CPI_M_PC_INTERNAL_27;
N_247 <= CPI_M_PC_INTERNAL_28;
N_248 <= CPI_M_PC_INTERNAL_29;
N_249 <= CPI_M_PC_INTERNAL_30;
N_250 <= CPI_M_INST_INTERNAL;
N_251 <= CPI_M_INST_INTERNAL_0;
N_252 <= CPI_M_INST_INTERNAL_1;
N_253 <= CPI_M_INST_INTERNAL_2;
N_254 <= CPI_M_INST_INTERNAL_3;
N_255 <= CPI_M_INST_INTERNAL_4;
N_256 <= CPI_M_INST_INTERNAL_5;
N_257 <= CPI_M_INST_INTERNAL_6;
N_258 <= CPI_M_INST_INTERNAL_7;
N_259 <= CPI_M_INST_INTERNAL_8;
N_260 <= CPI_M_INST_INTERNAL_9;
N_261 <= CPI_M_INST_INTERNAL_10;
N_262 <= CPI_M_INST_INTERNAL_11;
N_263 <= CPI_M_INST_INTERNAL_12;
N_264 <= CPI_M_INST_INTERNAL_13;
N_265 <= CPI_M_INST_INTERNAL_14;
N_266 <= CPI_M_INST_INTERNAL_15;
N_267 <= CPI_M_INST_INTERNAL_16;
N_268 <= CPI_M_INST_INTERNAL_17;
N_269 <= CPI_M_INST_INTERNAL_18;
N_270 <= CPI_M_INST_INTERNAL_19;
N_271 <= CPI_M_INST_INTERNAL_20;
N_272 <= CPI_M_INST_INTERNAL_21;
N_273 <= CPI_M_INST_INTERNAL_22;
N_274 <= CPI_M_INST_INTERNAL_23;
N_275 <= CPI_M_INST_INTERNAL_24;
N_276 <= CPI_M_INST_INTERNAL_25;
N_277 <= CPI_M_INST_INTERNAL_26;
N_278 <= CPI_M_INST_INTERNAL_27;
N_279 <= CPI_M_INST_INTERNAL_28;
N_280 <= CPI_M_INST_INTERNAL_29;
N_281 <= CPI_M_INST_INTERNAL_30;
N_282 <= CPI_M_CNT_INTERNAL;
N_283 <= CPI_M_CNT_INTERNAL_0;
N_284 <= CPI_M_TRAP_INTERNAL;
N_285 <= CPI_M_ANNUL_INTERNAL;
N_286 <= CPI_M_PV_INTERNAL;
N_287 <= CPI_X_PC_INTERNAL;
N_288 <= CPI_X_PC_INTERNAL_0;
N_289 <= CPI_X_PC_INTERNAL_1;
N_290 <= CPI_X_PC_INTERNAL_2;
N_291 <= CPI_X_PC_INTERNAL_3;
N_292 <= CPI_X_PC_INTERNAL_4;
N_293 <= CPI_X_PC_INTERNAL_5;
N_294 <= CPI_X_PC_INTERNAL_6;
N_295 <= CPI_X_PC_INTERNAL_7;
N_296 <= CPI_X_PC_INTERNAL_8;
N_297 <= CPI_X_PC_INTERNAL_9;
N_298 <= CPI_X_PC_INTERNAL_10;
N_299 <= CPI_X_PC_INTERNAL_11;
N_300 <= CPI_X_PC_INTERNAL_12;
N_301 <= CPI_X_PC_INTERNAL_13;
N_302 <= CPI_X_PC_INTERNAL_14;
N_303 <= CPI_X_PC_INTERNAL_15;
N_304 <= CPI_X_PC_INTERNAL_16;
N_305 <= CPI_X_PC_INTERNAL_17;
N_306 <= CPI_X_PC_INTERNAL_18;
N_307 <= CPI_X_PC_INTERNAL_19;
N_308 <= CPI_X_PC_INTERNAL_20;
N_309 <= CPI_X_PC_INTERNAL_21;
N_310 <= CPI_X_PC_INTERNAL_22;
N_311 <= CPI_X_PC_INTERNAL_23;
N_312 <= CPI_X_PC_INTERNAL_24;
N_313 <= CPI_X_PC_INTERNAL_25;
N_314 <= CPI_X_PC_INTERNAL_26;
N_315 <= CPI_X_PC_INTERNAL_27;
N_316 <= CPI_X_PC_INTERNAL_28;
N_317 <= CPI_X_PC_INTERNAL_29;
N_318 <= CPI_X_PC_INTERNAL_30;
N_319 <= CPI_X_INST_INTERNAL;
N_320 <= CPI_X_INST_INTERNAL_0;
N_321 <= CPI_X_INST_INTERNAL_1;
N_322 <= CPI_X_INST_INTERNAL_2;
N_323 <= CPI_X_INST_INTERNAL_3;
N_324 <= CPI_X_INST_INTERNAL_4;
N_325 <= CPI_X_INST_INTERNAL_5;
N_326 <= CPI_X_INST_INTERNAL_6;
N_327 <= CPI_X_INST_INTERNAL_7;
N_328 <= CPI_X_INST_INTERNAL_8;
N_329 <= CPI_X_INST_INTERNAL_9;
N_330 <= CPI_X_INST_INTERNAL_10;
N_331 <= CPI_X_INST_INTERNAL_11;
N_332 <= CPI_X_INST_INTERNAL_12;
N_333 <= CPI_X_INST_INTERNAL_13;
N_334 <= CPI_X_INST_INTERNAL_14;
N_335 <= CPI_X_INST_INTERNAL_15;
N_336 <= CPI_X_INST_INTERNAL_16;
N_337 <= CPI_X_INST_INTERNAL_17;
N_338 <= CPI_X_INST_INTERNAL_18;
N_339 <= CPI_X_INST_INTERNAL_19;
N_340 <= CPI_X_INST_INTERNAL_20;
N_341 <= CPI_X_INST_INTERNAL_21;
N_342 <= CPI_X_INST_INTERNAL_22;
N_343 <= CPI_X_INST_INTERNAL_23;
N_344 <= CPI_X_INST_INTERNAL_24;
N_345 <= CPI_X_INST_INTERNAL_25;
N_346 <= CPI_X_INST_INTERNAL_26;
N_347 <= CPI_X_INST_INTERNAL_27;
N_348 <= CPI_X_INST_INTERNAL_28;
N_349 <= CPI_X_INST_INTERNAL_29;
N_350 <= CPI_X_INST_INTERNAL_30;
N_351 <= CPI_X_CNT_INTERNAL;
N_352 <= CPI_X_CNT_INTERNAL_0;
N_353 <= CPI_X_TRAP_INTERNAL;
N_354 <= CPI_X_ANNUL_INTERNAL;
N_355 <= CPI_X_PV_INTERNAL;
N_356 <= CPI_LDDATA_INTERNAL;
N_357 <= CPI_LDDATA_INTERNAL_0;
N_358 <= CPI_LDDATA_INTERNAL_1;
N_359 <= CPI_LDDATA_INTERNAL_2;
N_360 <= CPI_LDDATA_INTERNAL_3;
N_361 <= CPI_LDDATA_INTERNAL_4;
N_362 <= CPI_LDDATA_INTERNAL_5;
N_363 <= CPI_LDDATA_INTERNAL_6;
N_364 <= CPI_LDDATA_INTERNAL_7;
N_365 <= CPI_LDDATA_INTERNAL_8;
N_366 <= CPI_LDDATA_INTERNAL_9;
N_367 <= CPI_LDDATA_INTERNAL_10;
N_368 <= CPI_LDDATA_INTERNAL_11;
N_369 <= CPI_LDDATA_INTERNAL_12;
N_370 <= CPI_LDDATA_INTERNAL_13;
N_371 <= CPI_LDDATA_INTERNAL_14;
N_372 <= CPI_LDDATA_INTERNAL_15;
N_373 <= CPI_LDDATA_INTERNAL_16;
N_374 <= CPI_LDDATA_INTERNAL_17;
N_375 <= CPI_LDDATA_INTERNAL_18;
N_376 <= CPI_LDDATA_INTERNAL_19;
N_377 <= CPI_LDDATA_INTERNAL_20;
N_378 <= CPI_LDDATA_INTERNAL_21;
N_379 <= CPI_LDDATA_INTERNAL_22;
N_380 <= CPI_LDDATA_INTERNAL_23;
N_381 <= CPI_LDDATA_INTERNAL_24;
N_382 <= CPI_LDDATA_INTERNAL_25;
N_383 <= CPI_LDDATA_INTERNAL_26;
N_384 <= CPI_LDDATA_INTERNAL_27;
N_385 <= CPI_LDDATA_INTERNAL_28;
N_386 <= CPI_LDDATA_INTERNAL_29;
N_387 <= CPI_LDDATA_INTERNAL_30;
N_388 <= CPI_DBG_ENABLE_INTERNAL;
N_389 <= CPI_DBG_WRITE_INTERNAL;
N_390 <= CPI_DBG_FSR_INTERNAL;
N_391 <= CPI_DBG_ADDR_INTERNAL;
N_392 <= CPI_DBG_ADDR_INTERNAL_0;
N_393 <= CPI_DBG_ADDR_INTERNAL_1;
N_394 <= CPI_DBG_ADDR_INTERNAL_2;
N_395 <= CPI_DBG_ADDR_INTERNAL_3;
N_396 <= CPI_DBG_DATA_INTERNAL;
N_397 <= CPI_DBG_DATA_INTERNAL_0;
N_398 <= CPI_DBG_DATA_INTERNAL_1;
N_399 <= CPI_DBG_DATA_INTERNAL_2;
N_400 <= CPI_DBG_DATA_INTERNAL_3;
N_401 <= CPI_DBG_DATA_INTERNAL_4;
N_402 <= CPI_DBG_DATA_INTERNAL_5;
N_403 <= CPI_DBG_DATA_INTERNAL_6;
N_404 <= CPI_DBG_DATA_INTERNAL_7;
N_405 <= CPI_DBG_DATA_INTERNAL_8;
N_406 <= CPI_DBG_DATA_INTERNAL_9;
N_407 <= CPI_DBG_DATA_INTERNAL_10;
N_408 <= CPI_DBG_DATA_INTERNAL_11;
N_409 <= CPI_DBG_DATA_INTERNAL_12;
N_410 <= CPI_DBG_DATA_INTERNAL_13;
N_411 <= CPI_DBG_DATA_INTERNAL_14;
N_412 <= CPI_DBG_DATA_INTERNAL_15;
N_413 <= CPI_DBG_DATA_INTERNAL_16;
N_414 <= CPI_DBG_DATA_INTERNAL_17;
N_415 <= CPI_DBG_DATA_INTERNAL_18;
N_416 <= CPI_DBG_DATA_INTERNAL_19;
N_417 <= CPI_DBG_DATA_INTERNAL_20;
N_418 <= CPI_DBG_DATA_INTERNAL_21;
N_419 <= CPI_DBG_DATA_INTERNAL_22;
N_420 <= CPI_DBG_DATA_INTERNAL_23;
N_421 <= CPI_DBG_DATA_INTERNAL_24;
N_422 <= CPI_DBG_DATA_INTERNAL_25;
N_423 <= CPI_DBG_DATA_INTERNAL_26;
N_424 <= CPI_DBG_DATA_INTERNAL_27;
N_425 <= CPI_DBG_DATA_INTERNAL_28;
N_426 <= CPI_DBG_DATA_INTERNAL_29;
N_427 <= CPI_DBG_DATA_INTERNAL_30;
N_0 <= CPO_DATAZ(0);
N_1_0 <= CPO_DATAZ(1);
N_2_0 <= CPO_DATAZ(2);
N_3_0 <= CPO_DATAZ(3);
N_4_0 <= CPO_DATAZ(4);
N_5_0 <= CPO_DATAZ(5);
N_6_0 <= CPO_DATAZ(6);
N_7_0 <= CPO_DATAZ(7);
N_8_0 <= CPO_DATAZ(8);
N_9_0 <= CPO_DATAZ(9);
N_10_0 <= CPO_DATAZ(10);
N_11_0 <= CPO_DATAZ(11);
N_12_0 <= CPO_DATAZ(12);
N_13_0 <= CPO_DATAZ(13);
N_14_0 <= CPO_DATAZ(14);
N_15_0 <= CPO_DATAZ(15);
N_16_0 <= CPO_DATAZ(16);
N_17_0 <= CPO_DATAZ(17);
N_18_0 <= CPO_DATAZ(18);
N_19_0 <= CPO_DATAZ(19);
N_20_0 <= CPO_DATAZ(20);
N_21_0 <= CPO_DATAZ(21);
N_22_0 <= CPO_DATAZ(22);
N_23_0 <= CPO_DATAZ(23);
N_24_0 <= CPO_DATAZ(24);
N_25_0 <= CPO_DATAZ(25);
N_26_0 <= CPO_DATAZ(26);
N_27_0 <= CPO_DATAZ(27);
N_28_0 <= CPO_DATAZ(28);
N_29_0 <= CPO_DATAZ(29);
N_30_0 <= CPO_DATAZ(30);
N_31_0 <= CPO_DATAZ(31);
N_32_0 <= CPO_EXCZ;
N_33_0 <= CPO_CCZ(0);
N_34_0 <= CPO_CCZ(1);
N_35_0 <= CPO_CCVZ;
N_36_0 <= CPO_LDLOCKZ;
N_37_0 <= CPO_HOLDNZ;
N_38_0 <= CPO_DBG_DATAZ(0);
N_39_0 <= CPO_DBG_DATAZ(1);
N_40_0 <= CPO_DBG_DATAZ(2);
N_41_0 <= CPO_DBG_DATAZ(3);
N_42_0 <= CPO_DBG_DATAZ(4);
N_43_0 <= CPO_DBG_DATAZ(5);
N_44_0 <= CPO_DBG_DATAZ(6);
N_45_0 <= CPO_DBG_DATAZ(7);
N_46_0 <= CPO_DBG_DATAZ(8);
N_47_0 <= CPO_DBG_DATAZ(9);
N_48_0 <= CPO_DBG_DATAZ(10);
N_49_0 <= CPO_DBG_DATAZ(11);
N_50_0 <= CPO_DBG_DATAZ(12);
N_51_0 <= CPO_DBG_DATAZ(13);
N_52_0 <= CPO_DBG_DATAZ(14);
N_53_0 <= CPO_DBG_DATAZ(15);
N_54_0 <= CPO_DBG_DATAZ(16);
N_55_0 <= CPO_DBG_DATAZ(17);
N_56_0 <= CPO_DBG_DATAZ(18);
N_57_0 <= CPO_DBG_DATAZ(19);
N_58_0 <= CPO_DBG_DATAZ(20);
N_59_0 <= CPO_DBG_DATAZ(21);
N_60_0 <= CPO_DBG_DATAZ(22);
N_61_0 <= CPO_DBG_DATAZ(23);
N_62_0 <= CPO_DBG_DATAZ(24);
N_63_0 <= CPO_DBG_DATAZ(25);
N_64_0 <= CPO_DBG_DATAZ(26);
N_65_0 <= CPO_DBG_DATAZ(27);
N_66_0 <= CPO_DBG_DATAZ(28);
N_67_0 <= CPO_DBG_DATAZ(29);
N_68_0 <= CPO_DBG_DATAZ(30);
N_69_0 <= CPO_DBG_DATAZ(31);
N_70_0 <= RFI2_RD1ADDRZ(0);
N_71_0 <= RFI2_RD1ADDRZ(1);
N_72_0 <= RFI2_RD1ADDRZ(2);
N_73_0 <= RFI2_RD1ADDRZ(3);
N_74_0 <= RFI2_RD2ADDRZ(0);
N_75_0 <= RFI2_RD2ADDRZ(1);
N_76_0 <= RFI2_RD2ADDRZ(2);
N_77_0 <= RFI2_RD2ADDRZ(3);
N_78_0 <= RFI2_WRADDRZ(0);
N_79_0 <= RFI2_WRADDRZ(1);
N_80_0 <= RFI2_WRADDRZ(2);
N_81_0 <= RFI2_WRADDRZ(3);
N_82_0 <= RFI1_WRDATAZ(0);
N_83_0 <= RFI1_WRDATAZ(1);
N_84_0 <= RFI1_WRDATAZ(2);
N_85_0 <= RFI1_WRDATAZ(3);
N_86_0 <= RFI1_WRDATAZ(4);
N_87_0 <= RFI1_WRDATAZ(5);
N_88_0 <= RFI1_WRDATAZ(6);
N_89_0 <= RFI1_WRDATAZ(7);
N_90_0 <= RFI1_WRDATAZ(8);
N_91_0 <= RFI1_WRDATAZ(9);
N_92_0 <= RFI1_WRDATAZ(10);
N_93_0 <= RFI1_WRDATAZ(11);
N_94_0 <= RFI1_WRDATAZ(12);
N_95_0 <= RFI1_WRDATAZ(13);
N_96_0 <= RFI1_WRDATAZ(14);
N_97_0 <= RFI1_WRDATAZ(15);
N_98_0 <= RFI1_WRDATAZ(16);
N_99_0 <= RFI1_WRDATAZ(17);
N_100_0 <= RFI1_WRDATAZ(18);
N_101_0 <= RFI1_WRDATAZ(19);
N_102_0 <= RFI1_WRDATAZ(20);
N_103_0 <= RFI1_WRDATAZ(21);
N_104_0 <= RFI1_WRDATAZ(22);
N_105_0 <= RFI1_WRDATAZ(23);
N_106_0 <= RFI1_WRDATAZ(24);
N_107_0 <= RFI1_WRDATAZ(25);
N_108_0 <= RFI1_WRDATAZ(26);
N_109_0 <= RFI1_WRDATAZ(27);
N_110_0 <= RFI1_WRDATAZ(28);
N_111_0 <= RFI1_WRDATAZ(29);
N_112_0 <= RFI1_WRDATAZ(30);
N_113_0 <= RFI1_WRDATAZ(31);
N_114_0 <= RFI1_REN1Z;
N_115_0 <= RFI1_REN2Z;
N_116_0 <= RFI1_WRENZ;
N_117_0 <= RFI2_RD1ADDRZ(0);
N_118_0 <= RFI2_RD1ADDRZ(1);
N_119_0 <= RFI2_RD1ADDRZ(2);
N_120_0 <= RFI2_RD1ADDRZ(3);
N_121_0 <= RFI2_RD2ADDRZ(0);
N_122_0 <= RFI2_RD2ADDRZ(1);
N_123_0 <= RFI2_RD2ADDRZ(2);
N_124_0 <= RFI2_RD2ADDRZ(3);
N_125_0 <= RFI2_WRADDRZ(0);
N_126_0 <= RFI2_WRADDRZ(1);
N_127_0 <= RFI2_WRADDRZ(2);
N_128_0 <= RFI2_WRADDRZ(3);
N_129_0 <= RFI2_WRDATAZ(0);
N_130_0 <= RFI2_WRDATAZ(1);
N_131_0 <= RFI2_WRDATAZ(2);
N_132_0 <= RFI2_WRDATAZ(3);
N_133_0 <= RFI2_WRDATAZ(4);
N_134_0 <= RFI2_WRDATAZ(5);
N_135_0 <= RFI2_WRDATAZ(6);
N_136_0 <= RFI2_WRDATAZ(7);
N_137_0 <= RFI2_WRDATAZ(8);
N_138_0 <= RFI2_WRDATAZ(9);
N_139_0 <= RFI2_WRDATAZ(10);
N_140_0 <= RFI2_WRDATAZ(11);
N_141_0 <= RFI2_WRDATAZ(12);
N_142_0 <= RFI2_WRDATAZ(13);
N_143_0 <= RFI2_WRDATAZ(14);
N_144_0 <= RFI2_WRDATAZ(15);
N_145_0 <= RFI2_WRDATAZ(16);
N_146_0 <= RFI2_WRDATAZ(17);
N_147_0 <= RFI2_WRDATAZ(18);
N_148_0 <= RFI2_WRDATAZ(19);
N_149_0 <= RFI2_WRDATAZ(20);
N_150_0 <= RFI2_WRDATAZ(21);
N_151_0 <= RFI2_WRDATAZ(22);
N_152_0 <= RFI2_WRDATAZ(23);
N_153_0 <= RFI2_WRDATAZ(24);
N_154_0 <= RFI2_WRDATAZ(25);
N_155_0 <= RFI2_WRDATAZ(26);
N_156_0 <= RFI2_WRDATAZ(27);
N_157_0 <= RFI2_WRDATAZ(28);
N_158_0 <= RFI2_WRDATAZ(29);
N_159_0 <= RFI2_WRDATAZ(30);
N_160_0 <= RFI2_WRDATAZ(31);
N_161_0 <= RFI2_REN1Z;
N_162_0 <= RFI2_REN2Z;
N_163_0 <= RFI2_WRENZ;
N_592 <= RFO1_DATA1_INTERNAL;
N_593 <= RFO1_DATA1_INTERNAL_0;
N_594 <= RFO1_DATA1_INTERNAL_1;
N_595 <= RFO1_DATA1_INTERNAL_2;
N_596 <= RFO1_DATA1_INTERNAL_3;
N_597 <= RFO1_DATA1_INTERNAL_4;
N_598 <= RFO1_DATA1_INTERNAL_5;
N_599 <= RFO1_DATA1_INTERNAL_6;
N_600 <= RFO1_DATA1_INTERNAL_7;
N_601 <= RFO1_DATA1_INTERNAL_8;
N_602 <= RFO1_DATA1_INTERNAL_9;
N_603 <= RFO1_DATA1_INTERNAL_10;
N_604 <= RFO1_DATA1_INTERNAL_11;
N_605 <= RFO1_DATA1_INTERNAL_12;
N_606 <= RFO1_DATA1_INTERNAL_13;
N_607 <= RFO1_DATA1_INTERNAL_14;
N_608 <= RFO1_DATA1_INTERNAL_15;
N_609 <= RFO1_DATA1_INTERNAL_16;
N_610 <= RFO1_DATA1_INTERNAL_17;
N_611 <= RFO1_DATA1_INTERNAL_18;
N_612 <= RFO1_DATA1_INTERNAL_19;
N_613 <= RFO1_DATA1_INTERNAL_20;
N_614 <= RFO1_DATA1_INTERNAL_21;
N_615 <= RFO1_DATA1_INTERNAL_22;
N_616 <= RFO1_DATA1_INTERNAL_23;
N_617 <= RFO1_DATA1_INTERNAL_24;
N_618 <= RFO1_DATA1_INTERNAL_25;
N_619 <= RFO1_DATA1_INTERNAL_26;
N_620 <= RFO1_DATA1_INTERNAL_27;
N_621 <= RFO1_DATA1_INTERNAL_28;
N_622 <= RFO1_DATA1_INTERNAL_29;
N_623 <= RFO1_DATA1_INTERNAL_30;
N_624 <= RFO1_DATA2_INTERNAL;
N_625 <= RFO1_DATA2_INTERNAL_0;
N_626 <= RFO1_DATA2_INTERNAL_1;
N_627 <= RFO1_DATA2_INTERNAL_2;
N_628 <= RFO1_DATA2_INTERNAL_3;
N_629 <= RFO1_DATA2_INTERNAL_4;
N_630 <= RFO1_DATA2_INTERNAL_5;
N_631 <= RFO1_DATA2_INTERNAL_6;
N_632 <= RFO1_DATA2_INTERNAL_7;
N_633 <= RFO1_DATA2_INTERNAL_8;
N_634 <= RFO1_DATA2_INTERNAL_9;
N_635 <= RFO1_DATA2_INTERNAL_10;
N_636 <= RFO1_DATA2_INTERNAL_11;
N_637 <= RFO1_DATA2_INTERNAL_12;
N_638 <= RFO1_DATA2_INTERNAL_13;
N_639 <= RFO1_DATA2_INTERNAL_14;
N_640 <= RFO1_DATA2_INTERNAL_15;
N_641 <= RFO1_DATA2_INTERNAL_16;
N_642 <= RFO1_DATA2_INTERNAL_17;
N_643 <= RFO1_DATA2_INTERNAL_18;
N_644 <= RFO1_DATA2_INTERNAL_19;
N_645 <= RFO1_DATA2_INTERNAL_20;
N_646 <= RFO1_DATA2_INTERNAL_21;
N_647 <= RFO1_DATA2_INTERNAL_22;
N_648 <= RFO1_DATA2_INTERNAL_23;
N_649 <= RFO1_DATA2_INTERNAL_24;
N_650 <= RFO1_DATA2_INTERNAL_25;
N_651 <= RFO1_DATA2_INTERNAL_26;
N_652 <= RFO1_DATA2_INTERNAL_27;
N_653 <= RFO1_DATA2_INTERNAL_28;
N_654 <= RFO1_DATA2_INTERNAL_29;
N_655 <= RFO1_DATA2_INTERNAL_30;
N_656 <= RFO2_DATA1_INTERNAL;
N_657 <= RFO2_DATA1_INTERNAL_0;
N_658 <= RFO2_DATA1_INTERNAL_1;
N_659 <= RFO2_DATA1_INTERNAL_2;
N_660 <= RFO2_DATA1_INTERNAL_3;
N_661 <= RFO2_DATA1_INTERNAL_4;
N_662 <= RFO2_DATA1_INTERNAL_5;
N_663 <= RFO2_DATA1_INTERNAL_6;
N_664 <= RFO2_DATA1_INTERNAL_7;
N_665 <= RFO2_DATA1_INTERNAL_8;
N_666 <= RFO2_DATA1_INTERNAL_9;
N_667 <= RFO2_DATA1_INTERNAL_10;
N_668 <= RFO2_DATA1_INTERNAL_11;
N_669 <= RFO2_DATA1_INTERNAL_12;
N_670 <= RFO2_DATA1_INTERNAL_13;
N_671 <= RFO2_DATA1_INTERNAL_14;
N_672 <= RFO2_DATA1_INTERNAL_15;
N_673 <= RFO2_DATA1_INTERNAL_16;
N_674 <= RFO2_DATA1_INTERNAL_17;
N_675 <= RFO2_DATA1_INTERNAL_18;
N_676 <= RFO2_DATA1_INTERNAL_19;
N_677 <= RFO2_DATA1_INTERNAL_20;
N_678 <= RFO2_DATA1_INTERNAL_21;
N_679 <= RFO2_DATA1_INTERNAL_22;
N_680 <= RFO2_DATA1_INTERNAL_23;
N_681 <= RFO2_DATA1_INTERNAL_24;
N_682 <= RFO2_DATA1_INTERNAL_25;
N_683 <= RFO2_DATA1_INTERNAL_26;
N_684 <= RFO2_DATA1_INTERNAL_27;
N_685 <= RFO2_DATA1_INTERNAL_28;
N_686 <= RFO2_DATA1_INTERNAL_29;
N_687 <= RFO2_DATA1_INTERNAL_30;
N_688 <= RFO2_DATA2_INTERNAL;
N_689 <= RFO2_DATA2_INTERNAL_0;
N_690 <= RFO2_DATA2_INTERNAL_1;
N_691 <= RFO2_DATA2_INTERNAL_2;
N_692 <= RFO2_DATA2_INTERNAL_3;
N_693 <= RFO2_DATA2_INTERNAL_4;
N_694 <= RFO2_DATA2_INTERNAL_5;
N_695 <= RFO2_DATA2_INTERNAL_6;
N_696 <= RFO2_DATA2_INTERNAL_7;
N_697 <= RFO2_DATA2_INTERNAL_8;
N_698 <= RFO2_DATA2_INTERNAL_9;
N_699 <= RFO2_DATA2_INTERNAL_10;
N_700 <= RFO2_DATA2_INTERNAL_11;
N_701 <= RFO2_DATA2_INTERNAL_12;
N_702 <= RFO2_DATA2_INTERNAL_13;
N_703 <= RFO2_DATA2_INTERNAL_14;
N_704 <= RFO2_DATA2_INTERNAL_15;
N_705 <= RFO2_DATA2_INTERNAL_16;
N_706 <= RFO2_DATA2_INTERNAL_17;
N_707 <= RFO2_DATA2_INTERNAL_18;
N_708 <= RFO2_DATA2_INTERNAL_19;
N_709 <= RFO2_DATA2_INTERNAL_20;
N_710 <= RFO2_DATA2_INTERNAL_21;
N_711 <= RFO2_DATA2_INTERNAL_22;
N_712 <= RFO2_DATA2_INTERNAL_23;
N_713 <= RFO2_DATA2_INTERNAL_24;
N_714 <= RFO2_DATA2_INTERNAL_25;
N_715 <= RFO2_DATA2_INTERNAL_26;
N_716 <= RFO2_DATA2_INTERNAL_27;
N_717 <= RFO2_DATA2_INTERNAL_28;
N_718 <= RFO2_DATA2_INTERNAL_29;
N_719 <= RFO2_DATA2_INTERNAL_30;
N_1_I <= not N_1;
\GRLFPC20.V.STATE_0_SQMUXA_1_X_I\ <= not \GRLFPC20.V.STATE_0_SQMUXA_1_X\;
\GRLFPC20.V.I.EXEC_0_SQMUXA_I\ <= not \GRLFPC20.V.I.EXEC_0_SQMUXA\;
\GRLFPC20.R.A.AFQ_I\ <= not \GRLFPC20.R.A.AFQ\;
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4_I\ <= not \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_1_SN_M4\;
\GRLFPC20.FPI.LDOP_I\ <= not \GRLFPC20.FPI.LDOP\;
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL_I\(78) <= not \GRLFPC20.GRFPUL_GEN0.GRLFPU0.R.PCTRL\(78);
\GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1_I\ <= not \GRLFPC20.GRFPUL_GEN0.GRLFPU0.RIN.DPATH_SN_M3_1\;
\GRLFPC20.COMB.UN2_HOLDN_I\ <= not \GRLFPC20.COMB.UN2_HOLDN\;
cpo_data(0) <= N_0;
cpo_data(1) <= N_1_0;
cpo_data(2) <= N_2_0;
cpo_data(3) <= N_3_0;
cpo_data(4) <= N_4_0;
cpo_data(5) <= N_5_0;
cpo_data(6) <= N_6_0;
cpo_data(7) <= N_7_0;
cpo_data(8) <= N_8_0;
cpo_data(9) <= N_9_0;
cpo_data(10) <= N_10_0;
cpo_data(11) <= N_11_0;
cpo_data(12) <= N_12_0;
cpo_data(13) <= N_13_0;
cpo_data(14) <= N_14_0;
cpo_data(15) <= N_15_0;
cpo_data(16) <= N_16_0;
cpo_data(17) <= N_17_0;
cpo_data(18) <= N_18_0;
cpo_data(19) <= N_19_0;
cpo_data(20) <= N_20_0;
cpo_data(21) <= N_21_0;
cpo_data(22) <= N_22_0;
cpo_data(23) <= N_23_0;
cpo_data(24) <= N_24_0;
cpo_data(25) <= N_25_0;
cpo_data(26) <= N_26_0;
cpo_data(27) <= N_27_0;
cpo_data(28) <= N_28_0;
cpo_data(29) <= N_29_0;
cpo_data(30) <= N_30_0;
cpo_data(31) <= N_31_0;
cpo_exc <= N_32_0;
cpo_cc(0) <= N_33_0;
cpo_cc(1) <= N_34_0;
cpo_ccv <= N_35_0;
cpo_ldlock <= N_36_0;
cpo_holdn <= N_37_0;
cpo_dbg_data(0) <= N_38_0;
cpo_dbg_data(1) <= N_39_0;
cpo_dbg_data(2) <= N_40_0;
cpo_dbg_data(3) <= N_41_0;
cpo_dbg_data(4) <= N_42_0;
cpo_dbg_data(5) <= N_43_0;
cpo_dbg_data(6) <= N_44_0;
cpo_dbg_data(7) <= N_45_0;
cpo_dbg_data(8) <= N_46_0;
cpo_dbg_data(9) <= N_47_0;
cpo_dbg_data(10) <= N_48_0;
cpo_dbg_data(11) <= N_49_0;
cpo_dbg_data(12) <= N_50_0;
cpo_dbg_data(13) <= N_51_0;
cpo_dbg_data(14) <= N_52_0;
cpo_dbg_data(15) <= N_53_0;
cpo_dbg_data(16) <= N_54_0;
cpo_dbg_data(17) <= N_55_0;
cpo_dbg_data(18) <= N_56_0;
cpo_dbg_data(19) <= N_57_0;
cpo_dbg_data(20) <= N_58_0;
cpo_dbg_data(21) <= N_59_0;
cpo_dbg_data(22) <= N_60_0;
cpo_dbg_data(23) <= N_61_0;
cpo_dbg_data(24) <= N_62_0;
cpo_dbg_data(25) <= N_63_0;
cpo_dbg_data(26) <= N_64_0;
cpo_dbg_data(27) <= N_65_0;
cpo_dbg_data(28) <= N_66_0;
cpo_dbg_data(29) <= N_67_0;
cpo_dbg_data(30) <= N_68_0;
cpo_dbg_data(31) <= N_69_0;
rfi1_rd1addr(0) <= N_70_0;
rfi1_rd1addr(1) <= N_71_0;
rfi1_rd1addr(2) <= N_72_0;
rfi1_rd1addr(3) <= N_73_0;
rfi1_rd2addr(0) <= N_74_0;
rfi1_rd2addr(1) <= N_75_0;
rfi1_rd2addr(2) <= N_76_0;
rfi1_rd2addr(3) <= N_77_0;
rfi1_wraddr(0) <= N_78_0;
rfi1_wraddr(1) <= N_79_0;
rfi1_wraddr(2) <= N_80_0;
rfi1_wraddr(3) <= N_81_0;
rfi1_wrdata(0) <= N_82_0;
rfi1_wrdata(1) <= N_83_0;
rfi1_wrdata(2) <= N_84_0;
rfi1_wrdata(3) <= N_85_0;
rfi1_wrdata(4) <= N_86_0;
rfi1_wrdata(5) <= N_87_0;
rfi1_wrdata(6) <= N_88_0;
rfi1_wrdata(7) <= N_89_0;
rfi1_wrdata(8) <= N_90_0;
rfi1_wrdata(9) <= N_91_0;
rfi1_wrdata(10) <= N_92_0;
rfi1_wrdata(11) <= N_93_0;
rfi1_wrdata(12) <= N_94_0;
rfi1_wrdata(13) <= N_95_0;
rfi1_wrdata(14) <= N_96_0;
rfi1_wrdata(15) <= N_97_0;
rfi1_wrdata(16) <= N_98_0;
rfi1_wrdata(17) <= N_99_0;
rfi1_wrdata(18) <= N_100_0;
rfi1_wrdata(19) <= N_101_0;
rfi1_wrdata(20) <= N_102_0;
rfi1_wrdata(21) <= N_103_0;
rfi1_wrdata(22) <= N_104_0;
rfi1_wrdata(23) <= N_105_0;
rfi1_wrdata(24) <= N_106_0;
rfi1_wrdata(25) <= N_107_0;
rfi1_wrdata(26) <= N_108_0;
rfi1_wrdata(27) <= N_109_0;
rfi1_wrdata(28) <= N_110_0;
rfi1_wrdata(29) <= N_111_0;
rfi1_wrdata(30) <= N_112_0;
rfi1_wrdata(31) <= N_113_0;
rfi1_ren1 <= N_114_0;
rfi1_ren2 <= N_115_0;
rfi1_wren <= N_116_0;
rfi2_rd1addr(0) <= N_117_0;
rfi2_rd1addr(1) <= N_118_0;
rfi2_rd1addr(2) <= N_119_0;
rfi2_rd1addr(3) <= N_120_0;
rfi2_rd2addr(0) <= N_121_0;
rfi2_rd2addr(1) <= N_122_0;
rfi2_rd2addr(2) <= N_123_0;
rfi2_rd2addr(3) <= N_124_0;
rfi2_wraddr(0) <= N_125_0;
rfi2_wraddr(1) <= N_126_0;
rfi2_wraddr(2) <= N_127_0;
rfi2_wraddr(3) <= N_128_0;
rfi2_wrdata(0) <= N_129_0;
rfi2_wrdata(1) <= N_130_0;
rfi2_wrdata(2) <= N_131_0;
rfi2_wrdata(3) <= N_132_0;
rfi2_wrdata(4) <= N_133_0;
rfi2_wrdata(5) <= N_134_0;
rfi2_wrdata(6) <= N_135_0;
rfi2_wrdata(7) <= N_136_0;
rfi2_wrdata(8) <= N_137_0;
rfi2_wrdata(9) <= N_138_0;
rfi2_wrdata(10) <= N_139_0;
rfi2_wrdata(11) <= N_140_0;
rfi2_wrdata(12) <= N_141_0;
rfi2_wrdata(13) <= N_142_0;
rfi2_wrdata(14) <= N_143_0;
rfi2_wrdata(15) <= N_144_0;
rfi2_wrdata(16) <= N_145_0;
rfi2_wrdata(17) <= N_146_0;
rfi2_wrdata(18) <= N_147_0;
rfi2_wrdata(19) <= N_148_0;
rfi2_wrdata(20) <= N_149_0;
rfi2_wrdata(21) <= N_150_0;
rfi2_wrdata(22) <= N_151_0;
rfi2_wrdata(23) <= N_152_0;
rfi2_wrdata(24) <= N_153_0;
rfi2_wrdata(25) <= N_154_0;
rfi2_wrdata(26) <= N_155_0;
rfi2_wrdata(27) <= N_156_0;
rfi2_wrdata(28) <= N_157_0;
rfi2_wrdata(29) <= N_158_0;
rfi2_wrdata(30) <= N_159_0;
rfi2_wrdata(31) <= N_160_0;
rfi2_ren1 <= N_161_0;
rfi2_ren2 <= N_162_0;
rfi2_wren <= N_163_0;
RST_INTERNAL <= rst;
CLK_INTERNAL <= clk;
HOLDN_INTERNAL <= holdn;
CPI_FLUSH_INTERNAL <= cpi_flush;
CPI_EXACK_INTERNAL <= cpi_exack;
CPI_A_RS1_INTERNAL <= cpi_a_rs1(0);
CPI_A_RS1_INTERNAL_0 <= cpi_a_rs1(1);
CPI_A_RS1_INTERNAL_1 <= cpi_a_rs1(2);
CPI_A_RS1_INTERNAL_2 <= cpi_a_rs1(3);
CPI_A_RS1_INTERNAL_3 <= cpi_a_rs1(4);
CPI_D_PC_INTERNAL <= cpi_d_pc(0);
CPI_D_PC_INTERNAL_0 <= cpi_d_pc(1);
CPI_D_PC_INTERNAL_1 <= cpi_d_pc(2);
CPI_D_PC_INTERNAL_2 <= cpi_d_pc(3);
CPI_D_PC_INTERNAL_3 <= cpi_d_pc(4);
CPI_D_PC_INTERNAL_4 <= cpi_d_pc(5);
CPI_D_PC_INTERNAL_5 <= cpi_d_pc(6);
CPI_D_PC_INTERNAL_6 <= cpi_d_pc(7);
CPI_D_PC_INTERNAL_7 <= cpi_d_pc(8);
CPI_D_PC_INTERNAL_8 <= cpi_d_pc(9);
CPI_D_PC_INTERNAL_9 <= cpi_d_pc(10);
CPI_D_PC_INTERNAL_10 <= cpi_d_pc(11);
CPI_D_PC_INTERNAL_11 <= cpi_d_pc(12);
CPI_D_PC_INTERNAL_12 <= cpi_d_pc(13);
CPI_D_PC_INTERNAL_13 <= cpi_d_pc(14);
CPI_D_PC_INTERNAL_14 <= cpi_d_pc(15);
CPI_D_PC_INTERNAL_15 <= cpi_d_pc(16);
CPI_D_PC_INTERNAL_16 <= cpi_d_pc(17);
CPI_D_PC_INTERNAL_17 <= cpi_d_pc(18);
CPI_D_PC_INTERNAL_18 <= cpi_d_pc(19);
CPI_D_PC_INTERNAL_19 <= cpi_d_pc(20);
CPI_D_PC_INTERNAL_20 <= cpi_d_pc(21);
CPI_D_PC_INTERNAL_21 <= cpi_d_pc(22);
CPI_D_PC_INTERNAL_22 <= cpi_d_pc(23);
CPI_D_PC_INTERNAL_23 <= cpi_d_pc(24);
CPI_D_PC_INTERNAL_24 <= cpi_d_pc(25);
CPI_D_PC_INTERNAL_25 <= cpi_d_pc(26);
CPI_D_PC_INTERNAL_26 <= cpi_d_pc(27);
CPI_D_PC_INTERNAL_27 <= cpi_d_pc(28);
CPI_D_PC_INTERNAL_28 <= cpi_d_pc(29);
CPI_D_PC_INTERNAL_29 <= cpi_d_pc(30);
CPI_D_PC_INTERNAL_30 <= cpi_d_pc(31);
CPI_D_INST_INTERNAL <= cpi_d_inst(0);
CPI_D_INST_INTERNAL_0 <= cpi_d_inst(1);
CPI_D_INST_INTERNAL_1 <= cpi_d_inst(2);
CPI_D_INST_INTERNAL_2 <= cpi_d_inst(3);
CPI_D_INST_INTERNAL_3 <= cpi_d_inst(4);
CPI_D_INST_INTERNAL_4 <= cpi_d_inst(5);
CPI_D_INST_INTERNAL_5 <= cpi_d_inst(6);
CPI_D_INST_INTERNAL_6 <= cpi_d_inst(7);
CPI_D_INST_INTERNAL_7 <= cpi_d_inst(8);
CPI_D_INST_INTERNAL_8 <= cpi_d_inst(9);
CPI_D_INST_INTERNAL_9 <= cpi_d_inst(10);
CPI_D_INST_INTERNAL_10 <= cpi_d_inst(11);
CPI_D_INST_INTERNAL_11 <= cpi_d_inst(12);
CPI_D_INST_INTERNAL_12 <= cpi_d_inst(13);
CPI_D_INST_INTERNAL_13 <= cpi_d_inst(14);
CPI_D_INST_INTERNAL_14 <= cpi_d_inst(15);
CPI_D_INST_INTERNAL_15 <= cpi_d_inst(16);
CPI_D_INST_INTERNAL_16 <= cpi_d_inst(17);
CPI_D_INST_INTERNAL_17 <= cpi_d_inst(18);
CPI_D_INST_INTERNAL_18 <= cpi_d_inst(19);
CPI_D_INST_INTERNAL_19 <= cpi_d_inst(20);
CPI_D_INST_INTERNAL_20 <= cpi_d_inst(21);
CPI_D_INST_INTERNAL_21 <= cpi_d_inst(22);
CPI_D_INST_INTERNAL_22 <= cpi_d_inst(23);
CPI_D_INST_INTERNAL_23 <= cpi_d_inst(24);
CPI_D_INST_INTERNAL_24 <= cpi_d_inst(25);
CPI_D_INST_INTERNAL_25 <= cpi_d_inst(26);
CPI_D_INST_INTERNAL_26 <= cpi_d_inst(27);
CPI_D_INST_INTERNAL_27 <= cpi_d_inst(28);
CPI_D_INST_INTERNAL_28 <= cpi_d_inst(29);
CPI_D_INST_INTERNAL_29 <= cpi_d_inst(30);
CPI_D_INST_INTERNAL_30 <= cpi_d_inst(31);
CPI_D_CNT_INTERNAL <= cpi_d_cnt(0);
CPI_D_CNT_INTERNAL_0 <= cpi_d_cnt(1);
CPI_D_TRAP_INTERNAL <= cpi_d_trap;
CPI_D_ANNUL_INTERNAL <= cpi_d_annul;
CPI_D_PV_INTERNAL <= cpi_d_pv;
CPI_A_PC_INTERNAL <= cpi_a_pc(0);
CPI_A_PC_INTERNAL_0 <= cpi_a_pc(1);
CPI_A_PC_INTERNAL_1 <= cpi_a_pc(2);
CPI_A_PC_INTERNAL_2 <= cpi_a_pc(3);
CPI_A_PC_INTERNAL_3 <= cpi_a_pc(4);
CPI_A_PC_INTERNAL_4 <= cpi_a_pc(5);
CPI_A_PC_INTERNAL_5 <= cpi_a_pc(6);
CPI_A_PC_INTERNAL_6 <= cpi_a_pc(7);
CPI_A_PC_INTERNAL_7 <= cpi_a_pc(8);
CPI_A_PC_INTERNAL_8 <= cpi_a_pc(9);
CPI_A_PC_INTERNAL_9 <= cpi_a_pc(10);
CPI_A_PC_INTERNAL_10 <= cpi_a_pc(11);
CPI_A_PC_INTERNAL_11 <= cpi_a_pc(12);
CPI_A_PC_INTERNAL_12 <= cpi_a_pc(13);
CPI_A_PC_INTERNAL_13 <= cpi_a_pc(14);
CPI_A_PC_INTERNAL_14 <= cpi_a_pc(15);
CPI_A_PC_INTERNAL_15 <= cpi_a_pc(16);
CPI_A_PC_INTERNAL_16 <= cpi_a_pc(17);
CPI_A_PC_INTERNAL_17 <= cpi_a_pc(18);
CPI_A_PC_INTERNAL_18 <= cpi_a_pc(19);
CPI_A_PC_INTERNAL_19 <= cpi_a_pc(20);
CPI_A_PC_INTERNAL_20 <= cpi_a_pc(21);
CPI_A_PC_INTERNAL_21 <= cpi_a_pc(22);
CPI_A_PC_INTERNAL_22 <= cpi_a_pc(23);
CPI_A_PC_INTERNAL_23 <= cpi_a_pc(24);
CPI_A_PC_INTERNAL_24 <= cpi_a_pc(25);
CPI_A_PC_INTERNAL_25 <= cpi_a_pc(26);
CPI_A_PC_INTERNAL_26 <= cpi_a_pc(27);
CPI_A_PC_INTERNAL_27 <= cpi_a_pc(28);
CPI_A_PC_INTERNAL_28 <= cpi_a_pc(29);
CPI_A_PC_INTERNAL_29 <= cpi_a_pc(30);
CPI_A_PC_INTERNAL_30 <= cpi_a_pc(31);
CPI_A_INST_INTERNAL <= cpi_a_inst(0);
CPI_A_INST_INTERNAL_0 <= cpi_a_inst(1);
CPI_A_INST_INTERNAL_1 <= cpi_a_inst(2);
CPI_A_INST_INTERNAL_2 <= cpi_a_inst(3);
CPI_A_INST_INTERNAL_3 <= cpi_a_inst(4);
CPI_A_INST_INTERNAL_4 <= cpi_a_inst(5);
CPI_A_INST_INTERNAL_5 <= cpi_a_inst(6);
CPI_A_INST_INTERNAL_6 <= cpi_a_inst(7);
CPI_A_INST_INTERNAL_7 <= cpi_a_inst(8);
CPI_A_INST_INTERNAL_8 <= cpi_a_inst(9);
CPI_A_INST_INTERNAL_9 <= cpi_a_inst(10);
CPI_A_INST_INTERNAL_10 <= cpi_a_inst(11);
CPI_A_INST_INTERNAL_11 <= cpi_a_inst(12);
CPI_A_INST_INTERNAL_12 <= cpi_a_inst(13);
CPI_A_INST_INTERNAL_13 <= cpi_a_inst(14);
CPI_A_INST_INTERNAL_14 <= cpi_a_inst(15);
CPI_A_INST_INTERNAL_15 <= cpi_a_inst(16);
CPI_A_INST_INTERNAL_16 <= cpi_a_inst(17);
CPI_A_INST_INTERNAL_17 <= cpi_a_inst(18);
CPI_A_INST_INTERNAL_18 <= cpi_a_inst(19);
CPI_A_INST_INTERNAL_19 <= cpi_a_inst(20);
CPI_A_INST_INTERNAL_20 <= cpi_a_inst(21);
CPI_A_INST_INTERNAL_21 <= cpi_a_inst(22);
CPI_A_INST_INTERNAL_22 <= cpi_a_inst(23);
CPI_A_INST_INTERNAL_23 <= cpi_a_inst(24);
CPI_A_INST_INTERNAL_24 <= cpi_a_inst(25);
CPI_A_INST_INTERNAL_25 <= cpi_a_inst(26);
CPI_A_INST_INTERNAL_26 <= cpi_a_inst(27);
CPI_A_INST_INTERNAL_27 <= cpi_a_inst(28);
CPI_A_INST_INTERNAL_28 <= cpi_a_inst(29);
CPI_A_INST_INTERNAL_29 <= cpi_a_inst(30);
CPI_A_INST_INTERNAL_30 <= cpi_a_inst(31);
CPI_A_CNT_INTERNAL <= cpi_a_cnt(0);
CPI_A_CNT_INTERNAL_0 <= cpi_a_cnt(1);
CPI_A_TRAP_INTERNAL <= cpi_a_trap;
CPI_A_ANNUL_INTERNAL <= cpi_a_annul;
CPI_A_PV_INTERNAL <= cpi_a_pv;
CPI_E_PC_INTERNAL <= cpi_e_pc(0);
CPI_E_PC_INTERNAL_0 <= cpi_e_pc(1);
CPI_E_PC_INTERNAL_1 <= cpi_e_pc(2);
CPI_E_PC_INTERNAL_2 <= cpi_e_pc(3);
CPI_E_PC_INTERNAL_3 <= cpi_e_pc(4);
CPI_E_PC_INTERNAL_4 <= cpi_e_pc(5);
CPI_E_PC_INTERNAL_5 <= cpi_e_pc(6);
CPI_E_PC_INTERNAL_6 <= cpi_e_pc(7);
CPI_E_PC_INTERNAL_7 <= cpi_e_pc(8);
CPI_E_PC_INTERNAL_8 <= cpi_e_pc(9);
CPI_E_PC_INTERNAL_9 <= cpi_e_pc(10);
CPI_E_PC_INTERNAL_10 <= cpi_e_pc(11);
CPI_E_PC_INTERNAL_11 <= cpi_e_pc(12);
CPI_E_PC_INTERNAL_12 <= cpi_e_pc(13);
CPI_E_PC_INTERNAL_13 <= cpi_e_pc(14);
CPI_E_PC_INTERNAL_14 <= cpi_e_pc(15);
CPI_E_PC_INTERNAL_15 <= cpi_e_pc(16);
CPI_E_PC_INTERNAL_16 <= cpi_e_pc(17);
CPI_E_PC_INTERNAL_17 <= cpi_e_pc(18);
CPI_E_PC_INTERNAL_18 <= cpi_e_pc(19);
CPI_E_PC_INTERNAL_19 <= cpi_e_pc(20);
CPI_E_PC_INTERNAL_20 <= cpi_e_pc(21);
CPI_E_PC_INTERNAL_21 <= cpi_e_pc(22);
CPI_E_PC_INTERNAL_22 <= cpi_e_pc(23);
CPI_E_PC_INTERNAL_23 <= cpi_e_pc(24);
CPI_E_PC_INTERNAL_24 <= cpi_e_pc(25);
CPI_E_PC_INTERNAL_25 <= cpi_e_pc(26);
CPI_E_PC_INTERNAL_26 <= cpi_e_pc(27);
CPI_E_PC_INTERNAL_27 <= cpi_e_pc(28);
CPI_E_PC_INTERNAL_28 <= cpi_e_pc(29);
CPI_E_PC_INTERNAL_29 <= cpi_e_pc(30);
CPI_E_PC_INTERNAL_30 <= cpi_e_pc(31);
CPI_E_INST_INTERNAL <= cpi_e_inst(0);
CPI_E_INST_INTERNAL_0 <= cpi_e_inst(1);
CPI_E_INST_INTERNAL_1 <= cpi_e_inst(2);
CPI_E_INST_INTERNAL_2 <= cpi_e_inst(3);
CPI_E_INST_INTERNAL_3 <= cpi_e_inst(4);
CPI_E_INST_INTERNAL_4 <= cpi_e_inst(5);
CPI_E_INST_INTERNAL_5 <= cpi_e_inst(6);
CPI_E_INST_INTERNAL_6 <= cpi_e_inst(7);
CPI_E_INST_INTERNAL_7 <= cpi_e_inst(8);
CPI_E_INST_INTERNAL_8 <= cpi_e_inst(9);
CPI_E_INST_INTERNAL_9 <= cpi_e_inst(10);
CPI_E_INST_INTERNAL_10 <= cpi_e_inst(11);
CPI_E_INST_INTERNAL_11 <= cpi_e_inst(12);
CPI_E_INST_INTERNAL_12 <= cpi_e_inst(13);
CPI_E_INST_INTERNAL_13 <= cpi_e_inst(14);
CPI_E_INST_INTERNAL_14 <= cpi_e_inst(15);
CPI_E_INST_INTERNAL_15 <= cpi_e_inst(16);
CPI_E_INST_INTERNAL_16 <= cpi_e_inst(17);
CPI_E_INST_INTERNAL_17 <= cpi_e_inst(18);
CPI_E_INST_INTERNAL_18 <= cpi_e_inst(19);
CPI_E_INST_INTERNAL_19 <= cpi_e_inst(20);
CPI_E_INST_INTERNAL_20 <= cpi_e_inst(21);
CPI_E_INST_INTERNAL_21 <= cpi_e_inst(22);
CPI_E_INST_INTERNAL_22 <= cpi_e_inst(23);
CPI_E_INST_INTERNAL_23 <= cpi_e_inst(24);
CPI_E_INST_INTERNAL_24 <= cpi_e_inst(25);
CPI_E_INST_INTERNAL_25 <= cpi_e_inst(26);
CPI_E_INST_INTERNAL_26 <= cpi_e_inst(27);
CPI_E_INST_INTERNAL_27 <= cpi_e_inst(28);
CPI_E_INST_INTERNAL_28 <= cpi_e_inst(29);
CPI_E_INST_INTERNAL_29 <= cpi_e_inst(30);
CPI_E_INST_INTERNAL_30 <= cpi_e_inst(31);
CPI_E_CNT_INTERNAL <= cpi_e_cnt(0);
CPI_E_CNT_INTERNAL_0 <= cpi_e_cnt(1);
CPI_E_TRAP_INTERNAL <= cpi_e_trap;
CPI_E_ANNUL_INTERNAL <= cpi_e_annul;
CPI_E_PV_INTERNAL <= cpi_e_pv;
CPI_M_PC_INTERNAL <= cpi_m_pc(0);
CPI_M_PC_INTERNAL_0 <= cpi_m_pc(1);
CPI_M_PC_INTERNAL_1 <= cpi_m_pc(2);
CPI_M_PC_INTERNAL_2 <= cpi_m_pc(3);
CPI_M_PC_INTERNAL_3 <= cpi_m_pc(4);
CPI_M_PC_INTERNAL_4 <= cpi_m_pc(5);
CPI_M_PC_INTERNAL_5 <= cpi_m_pc(6);
CPI_M_PC_INTERNAL_6 <= cpi_m_pc(7);
CPI_M_PC_INTERNAL_7 <= cpi_m_pc(8);
CPI_M_PC_INTERNAL_8 <= cpi_m_pc(9);
CPI_M_PC_INTERNAL_9 <= cpi_m_pc(10);
CPI_M_PC_INTERNAL_10 <= cpi_m_pc(11);
CPI_M_PC_INTERNAL_11 <= cpi_m_pc(12);
CPI_M_PC_INTERNAL_12 <= cpi_m_pc(13);
CPI_M_PC_INTERNAL_13 <= cpi_m_pc(14);
CPI_M_PC_INTERNAL_14 <= cpi_m_pc(15);
CPI_M_PC_INTERNAL_15 <= cpi_m_pc(16);
CPI_M_PC_INTERNAL_16 <= cpi_m_pc(17);
CPI_M_PC_INTERNAL_17 <= cpi_m_pc(18);
CPI_M_PC_INTERNAL_18 <= cpi_m_pc(19);
CPI_M_PC_INTERNAL_19 <= cpi_m_pc(20);
CPI_M_PC_INTERNAL_20 <= cpi_m_pc(21);
CPI_M_PC_INTERNAL_21 <= cpi_m_pc(22);
CPI_M_PC_INTERNAL_22 <= cpi_m_pc(23);
CPI_M_PC_INTERNAL_23 <= cpi_m_pc(24);
CPI_M_PC_INTERNAL_24 <= cpi_m_pc(25);
CPI_M_PC_INTERNAL_25 <= cpi_m_pc(26);
CPI_M_PC_INTERNAL_26 <= cpi_m_pc(27);
CPI_M_PC_INTERNAL_27 <= cpi_m_pc(28);
CPI_M_PC_INTERNAL_28 <= cpi_m_pc(29);
CPI_M_PC_INTERNAL_29 <= cpi_m_pc(30);
CPI_M_PC_INTERNAL_30 <= cpi_m_pc(31);
CPI_M_INST_INTERNAL <= cpi_m_inst(0);
CPI_M_INST_INTERNAL_0 <= cpi_m_inst(1);
CPI_M_INST_INTERNAL_1 <= cpi_m_inst(2);
CPI_M_INST_INTERNAL_2 <= cpi_m_inst(3);
CPI_M_INST_INTERNAL_3 <= cpi_m_inst(4);
CPI_M_INST_INTERNAL_4 <= cpi_m_inst(5);
CPI_M_INST_INTERNAL_5 <= cpi_m_inst(6);
CPI_M_INST_INTERNAL_6 <= cpi_m_inst(7);
CPI_M_INST_INTERNAL_7 <= cpi_m_inst(8);
CPI_M_INST_INTERNAL_8 <= cpi_m_inst(9);
CPI_M_INST_INTERNAL_9 <= cpi_m_inst(10);
CPI_M_INST_INTERNAL_10 <= cpi_m_inst(11);
CPI_M_INST_INTERNAL_11 <= cpi_m_inst(12);
CPI_M_INST_INTERNAL_12 <= cpi_m_inst(13);
CPI_M_INST_INTERNAL_13 <= cpi_m_inst(14);
CPI_M_INST_INTERNAL_14 <= cpi_m_inst(15);
CPI_M_INST_INTERNAL_15 <= cpi_m_inst(16);
CPI_M_INST_INTERNAL_16 <= cpi_m_inst(17);
CPI_M_INST_INTERNAL_17 <= cpi_m_inst(18);
CPI_M_INST_INTERNAL_18 <= cpi_m_inst(19);
CPI_M_INST_INTERNAL_19 <= cpi_m_inst(20);
CPI_M_INST_INTERNAL_20 <= cpi_m_inst(21);
CPI_M_INST_INTERNAL_21 <= cpi_m_inst(22);
CPI_M_INST_INTERNAL_22 <= cpi_m_inst(23);
CPI_M_INST_INTERNAL_23 <= cpi_m_inst(24);
CPI_M_INST_INTERNAL_24 <= cpi_m_inst(25);
CPI_M_INST_INTERNAL_25 <= cpi_m_inst(26);
CPI_M_INST_INTERNAL_26 <= cpi_m_inst(27);
CPI_M_INST_INTERNAL_27 <= cpi_m_inst(28);
CPI_M_INST_INTERNAL_28 <= cpi_m_inst(29);
CPI_M_INST_INTERNAL_29 <= cpi_m_inst(30);
CPI_M_INST_INTERNAL_30 <= cpi_m_inst(31);
CPI_M_CNT_INTERNAL <= cpi_m_cnt(0);
CPI_M_CNT_INTERNAL_0 <= cpi_m_cnt(1);
CPI_M_TRAP_INTERNAL <= cpi_m_trap;
CPI_M_ANNUL_INTERNAL <= cpi_m_annul;
CPI_M_PV_INTERNAL <= cpi_m_pv;
CPI_X_PC_INTERNAL <= cpi_x_pc(0);
CPI_X_PC_INTERNAL_0 <= cpi_x_pc(1);
CPI_X_PC_INTERNAL_1 <= cpi_x_pc(2);
CPI_X_PC_INTERNAL_2 <= cpi_x_pc(3);
CPI_X_PC_INTERNAL_3 <= cpi_x_pc(4);
CPI_X_PC_INTERNAL_4 <= cpi_x_pc(5);
CPI_X_PC_INTERNAL_5 <= cpi_x_pc(6);
CPI_X_PC_INTERNAL_6 <= cpi_x_pc(7);
CPI_X_PC_INTERNAL_7 <= cpi_x_pc(8);
CPI_X_PC_INTERNAL_8 <= cpi_x_pc(9);
CPI_X_PC_INTERNAL_9 <= cpi_x_pc(10);
CPI_X_PC_INTERNAL_10 <= cpi_x_pc(11);
CPI_X_PC_INTERNAL_11 <= cpi_x_pc(12);
CPI_X_PC_INTERNAL_12 <= cpi_x_pc(13);
CPI_X_PC_INTERNAL_13 <= cpi_x_pc(14);
CPI_X_PC_INTERNAL_14 <= cpi_x_pc(15);
CPI_X_PC_INTERNAL_15 <= cpi_x_pc(16);
CPI_X_PC_INTERNAL_16 <= cpi_x_pc(17);
CPI_X_PC_INTERNAL_17 <= cpi_x_pc(18);
CPI_X_PC_INTERNAL_18 <= cpi_x_pc(19);
CPI_X_PC_INTERNAL_19 <= cpi_x_pc(20);
CPI_X_PC_INTERNAL_20 <= cpi_x_pc(21);
CPI_X_PC_INTERNAL_21 <= cpi_x_pc(22);
CPI_X_PC_INTERNAL_22 <= cpi_x_pc(23);
CPI_X_PC_INTERNAL_23 <= cpi_x_pc(24);
CPI_X_PC_INTERNAL_24 <= cpi_x_pc(25);
CPI_X_PC_INTERNAL_25 <= cpi_x_pc(26);
CPI_X_PC_INTERNAL_26 <= cpi_x_pc(27);
CPI_X_PC_INTERNAL_27 <= cpi_x_pc(28);
CPI_X_PC_INTERNAL_28 <= cpi_x_pc(29);
CPI_X_PC_INTERNAL_29 <= cpi_x_pc(30);
CPI_X_PC_INTERNAL_30 <= cpi_x_pc(31);
CPI_X_INST_INTERNAL <= cpi_x_inst(0);
CPI_X_INST_INTERNAL_0 <= cpi_x_inst(1);
CPI_X_INST_INTERNAL_1 <= cpi_x_inst(2);
CPI_X_INST_INTERNAL_2 <= cpi_x_inst(3);
CPI_X_INST_INTERNAL_3 <= cpi_x_inst(4);
CPI_X_INST_INTERNAL_4 <= cpi_x_inst(5);
CPI_X_INST_INTERNAL_5 <= cpi_x_inst(6);
CPI_X_INST_INTERNAL_6 <= cpi_x_inst(7);
CPI_X_INST_INTERNAL_7 <= cpi_x_inst(8);
CPI_X_INST_INTERNAL_8 <= cpi_x_inst(9);
CPI_X_INST_INTERNAL_9 <= cpi_x_inst(10);
CPI_X_INST_INTERNAL_10 <= cpi_x_inst(11);
CPI_X_INST_INTERNAL_11 <= cpi_x_inst(12);
CPI_X_INST_INTERNAL_12 <= cpi_x_inst(13);
CPI_X_INST_INTERNAL_13 <= cpi_x_inst(14);
CPI_X_INST_INTERNAL_14 <= cpi_x_inst(15);
CPI_X_INST_INTERNAL_15 <= cpi_x_inst(16);
CPI_X_INST_INTERNAL_16 <= cpi_x_inst(17);
CPI_X_INST_INTERNAL_17 <= cpi_x_inst(18);
CPI_X_INST_INTERNAL_18 <= cpi_x_inst(19);
CPI_X_INST_INTERNAL_19 <= cpi_x_inst(20);
CPI_X_INST_INTERNAL_20 <= cpi_x_inst(21);
CPI_X_INST_INTERNAL_21 <= cpi_x_inst(22);
CPI_X_INST_INTERNAL_22 <= cpi_x_inst(23);
CPI_X_INST_INTERNAL_23 <= cpi_x_inst(24);
CPI_X_INST_INTERNAL_24 <= cpi_x_inst(25);
CPI_X_INST_INTERNAL_25 <= cpi_x_inst(26);
CPI_X_INST_INTERNAL_26 <= cpi_x_inst(27);
CPI_X_INST_INTERNAL_27 <= cpi_x_inst(28);
CPI_X_INST_INTERNAL_28 <= cpi_x_inst(29);
CPI_X_INST_INTERNAL_29 <= cpi_x_inst(30);
CPI_X_INST_INTERNAL_30 <= cpi_x_inst(31);
CPI_X_CNT_INTERNAL <= cpi_x_cnt(0);
CPI_X_CNT_INTERNAL_0 <= cpi_x_cnt(1);
CPI_X_TRAP_INTERNAL <= cpi_x_trap;
CPI_X_ANNUL_INTERNAL <= cpi_x_annul;
CPI_X_PV_INTERNAL <= cpi_x_pv;
CPI_LDDATA_INTERNAL <= cpi_lddata(0);
CPI_LDDATA_INTERNAL_0 <= cpi_lddata(1);
CPI_LDDATA_INTERNAL_1 <= cpi_lddata(2);
CPI_LDDATA_INTERNAL_2 <= cpi_lddata(3);
CPI_LDDATA_INTERNAL_3 <= cpi_lddata(4);
CPI_LDDATA_INTERNAL_4 <= cpi_lddata(5);
CPI_LDDATA_INTERNAL_5 <= cpi_lddata(6);
CPI_LDDATA_INTERNAL_6 <= cpi_lddata(7);
CPI_LDDATA_INTERNAL_7 <= cpi_lddata(8);
CPI_LDDATA_INTERNAL_8 <= cpi_lddata(9);
CPI_LDDATA_INTERNAL_9 <= cpi_lddata(10);
CPI_LDDATA_INTERNAL_10 <= cpi_lddata(11);
CPI_LDDATA_INTERNAL_11 <= cpi_lddata(12);
CPI_LDDATA_INTERNAL_12 <= cpi_lddata(13);
CPI_LDDATA_INTERNAL_13 <= cpi_lddata(14);
CPI_LDDATA_INTERNAL_14 <= cpi_lddata(15);
CPI_LDDATA_INTERNAL_15 <= cpi_lddata(16);
CPI_LDDATA_INTERNAL_16 <= cpi_lddata(17);
CPI_LDDATA_INTERNAL_17 <= cpi_lddata(18);
CPI_LDDATA_INTERNAL_18 <= cpi_lddata(19);
CPI_LDDATA_INTERNAL_19 <= cpi_lddata(20);
CPI_LDDATA_INTERNAL_20 <= cpi_lddata(21);
CPI_LDDATA_INTERNAL_21 <= cpi_lddata(22);
CPI_LDDATA_INTERNAL_22 <= cpi_lddata(23);
CPI_LDDATA_INTERNAL_23 <= cpi_lddata(24);
CPI_LDDATA_INTERNAL_24 <= cpi_lddata(25);
CPI_LDDATA_INTERNAL_25 <= cpi_lddata(26);
CPI_LDDATA_INTERNAL_26 <= cpi_lddata(27);
CPI_LDDATA_INTERNAL_27 <= cpi_lddata(28);
CPI_LDDATA_INTERNAL_28 <= cpi_lddata(29);
CPI_LDDATA_INTERNAL_29 <= cpi_lddata(30);
CPI_LDDATA_INTERNAL_30 <= cpi_lddata(31);
CPI_DBG_ENABLE_INTERNAL <= cpi_dbg_enable;
CPI_DBG_WRITE_INTERNAL <= cpi_dbg_write;
CPI_DBG_FSR_INTERNAL <= cpi_dbg_fsr;
CPI_DBG_ADDR_INTERNAL <= cpi_dbg_addr(0);
CPI_DBG_ADDR_INTERNAL_0 <= cpi_dbg_addr(1);
CPI_DBG_ADDR_INTERNAL_1 <= cpi_dbg_addr(2);
CPI_DBG_ADDR_INTERNAL_2 <= cpi_dbg_addr(3);
CPI_DBG_ADDR_INTERNAL_3 <= cpi_dbg_addr(4);
CPI_DBG_DATA_INTERNAL <= cpi_dbg_data(0);
CPI_DBG_DATA_INTERNAL_0 <= cpi_dbg_data(1);
CPI_DBG_DATA_INTERNAL_1 <= cpi_dbg_data(2);
CPI_DBG_DATA_INTERNAL_2 <= cpi_dbg_data(3);
CPI_DBG_DATA_INTERNAL_3 <= cpi_dbg_data(4);
CPI_DBG_DATA_INTERNAL_4 <= cpi_dbg_data(5);
CPI_DBG_DATA_INTERNAL_5 <= cpi_dbg_data(6);
CPI_DBG_DATA_INTERNAL_6 <= cpi_dbg_data(7);
CPI_DBG_DATA_INTERNAL_7 <= cpi_dbg_data(8);
CPI_DBG_DATA_INTERNAL_8 <= cpi_dbg_data(9);
CPI_DBG_DATA_INTERNAL_9 <= cpi_dbg_data(10);
CPI_DBG_DATA_INTERNAL_10 <= cpi_dbg_data(11);
CPI_DBG_DATA_INTERNAL_11 <= cpi_dbg_data(12);
CPI_DBG_DATA_INTERNAL_12 <= cpi_dbg_data(13);
CPI_DBG_DATA_INTERNAL_13 <= cpi_dbg_data(14);
CPI_DBG_DATA_INTERNAL_14 <= cpi_dbg_data(15);
CPI_DBG_DATA_INTERNAL_15 <= cpi_dbg_data(16);
CPI_DBG_DATA_INTERNAL_16 <= cpi_dbg_data(17);
CPI_DBG_DATA_INTERNAL_17 <= cpi_dbg_data(18);
CPI_DBG_DATA_INTERNAL_18 <= cpi_dbg_data(19);
CPI_DBG_DATA_INTERNAL_19 <= cpi_dbg_data(20);
CPI_DBG_DATA_INTERNAL_20 <= cpi_dbg_data(21);
CPI_DBG_DATA_INTERNAL_21 <= cpi_dbg_data(22);
CPI_DBG_DATA_INTERNAL_22 <= cpi_dbg_data(23);
CPI_DBG_DATA_INTERNAL_23 <= cpi_dbg_data(24);
CPI_DBG_DATA_INTERNAL_24 <= cpi_dbg_data(25);
CPI_DBG_DATA_INTERNAL_25 <= cpi_dbg_data(26);
CPI_DBG_DATA_INTERNAL_26 <= cpi_dbg_data(27);
CPI_DBG_DATA_INTERNAL_27 <= cpi_dbg_data(28);
CPI_DBG_DATA_INTERNAL_28 <= cpi_dbg_data(29);
CPI_DBG_DATA_INTERNAL_29 <= cpi_dbg_data(30);
CPI_DBG_DATA_INTERNAL_30 <= cpi_dbg_data(31);
RFO1_DATA1_INTERNAL <= rfo1_data1(0);
RFO1_DATA1_INTERNAL_0 <= rfo1_data1(1);
RFO1_DATA1_INTERNAL_1 <= rfo1_data1(2);
RFO1_DATA1_INTERNAL_2 <= rfo1_data1(3);
RFO1_DATA1_INTERNAL_3 <= rfo1_data1(4);
RFO1_DATA1_INTERNAL_4 <= rfo1_data1(5);
RFO1_DATA1_INTERNAL_5 <= rfo1_data1(6);
RFO1_DATA1_INTERNAL_6 <= rfo1_data1(7);
RFO1_DATA1_INTERNAL_7 <= rfo1_data1(8);
RFO1_DATA1_INTERNAL_8 <= rfo1_data1(9);
RFO1_DATA1_INTERNAL_9 <= rfo1_data1(10);
RFO1_DATA1_INTERNAL_10 <= rfo1_data1(11);
RFO1_DATA1_INTERNAL_11 <= rfo1_data1(12);
RFO1_DATA1_INTERNAL_12 <= rfo1_data1(13);
RFO1_DATA1_INTERNAL_13 <= rfo1_data1(14);
RFO1_DATA1_INTERNAL_14 <= rfo1_data1(15);
RFO1_DATA1_INTERNAL_15 <= rfo1_data1(16);
RFO1_DATA1_INTERNAL_16 <= rfo1_data1(17);
RFO1_DATA1_INTERNAL_17 <= rfo1_data1(18);
RFO1_DATA1_INTERNAL_18 <= rfo1_data1(19);
RFO1_DATA1_INTERNAL_19 <= rfo1_data1(20);
RFO1_DATA1_INTERNAL_20 <= rfo1_data1(21);
RFO1_DATA1_INTERNAL_21 <= rfo1_data1(22);
RFO1_DATA1_INTERNAL_22 <= rfo1_data1(23);
RFO1_DATA1_INTERNAL_23 <= rfo1_data1(24);
RFO1_DATA1_INTERNAL_24 <= rfo1_data1(25);
RFO1_DATA1_INTERNAL_25 <= rfo1_data1(26);
RFO1_DATA1_INTERNAL_26 <= rfo1_data1(27);
RFO1_DATA1_INTERNAL_27 <= rfo1_data1(28);
RFO1_DATA1_INTERNAL_28 <= rfo1_data1(29);
RFO1_DATA1_INTERNAL_29 <= rfo1_data1(30);
RFO1_DATA1_INTERNAL_30 <= rfo1_data1(31);
RFO1_DATA2_INTERNAL <= rfo1_data2(0);
RFO1_DATA2_INTERNAL_0 <= rfo1_data2(1);
RFO1_DATA2_INTERNAL_1 <= rfo1_data2(2);
RFO1_DATA2_INTERNAL_2 <= rfo1_data2(3);
RFO1_DATA2_INTERNAL_3 <= rfo1_data2(4);
RFO1_DATA2_INTERNAL_4 <= rfo1_data2(5);
RFO1_DATA2_INTERNAL_5 <= rfo1_data2(6);
RFO1_DATA2_INTERNAL_6 <= rfo1_data2(7);
RFO1_DATA2_INTERNAL_7 <= rfo1_data2(8);
RFO1_DATA2_INTERNAL_8 <= rfo1_data2(9);
RFO1_DATA2_INTERNAL_9 <= rfo1_data2(10);
RFO1_DATA2_INTERNAL_10 <= rfo1_data2(11);
RFO1_DATA2_INTERNAL_11 <= rfo1_data2(12);
RFO1_DATA2_INTERNAL_12 <= rfo1_data2(13);
RFO1_DATA2_INTERNAL_13 <= rfo1_data2(14);
RFO1_DATA2_INTERNAL_14 <= rfo1_data2(15);
RFO1_DATA2_INTERNAL_15 <= rfo1_data2(16);
RFO1_DATA2_INTERNAL_16 <= rfo1_data2(17);
RFO1_DATA2_INTERNAL_17 <= rfo1_data2(18);
RFO1_DATA2_INTERNAL_18 <= rfo1_data2(19);
RFO1_DATA2_INTERNAL_19 <= rfo1_data2(20);
RFO1_DATA2_INTERNAL_20 <= rfo1_data2(21);
RFO1_DATA2_INTERNAL_21 <= rfo1_data2(22);
RFO1_DATA2_INTERNAL_22 <= rfo1_data2(23);
RFO1_DATA2_INTERNAL_23 <= rfo1_data2(24);
RFO1_DATA2_INTERNAL_24 <= rfo1_data2(25);
RFO1_DATA2_INTERNAL_25 <= rfo1_data2(26);
RFO1_DATA2_INTERNAL_26 <= rfo1_data2(27);
RFO1_DATA2_INTERNAL_27 <= rfo1_data2(28);
RFO1_DATA2_INTERNAL_28 <= rfo1_data2(29);
RFO1_DATA2_INTERNAL_29 <= rfo1_data2(30);
RFO1_DATA2_INTERNAL_30 <= rfo1_data2(31);
RFO2_DATA1_INTERNAL <= rfo2_data1(0);
RFO2_DATA1_INTERNAL_0 <= rfo2_data1(1);
RFO2_DATA1_INTERNAL_1 <= rfo2_data1(2);
RFO2_DATA1_INTERNAL_2 <= rfo2_data1(3);
RFO2_DATA1_INTERNAL_3 <= rfo2_data1(4);
RFO2_DATA1_INTERNAL_4 <= rfo2_data1(5);
RFO2_DATA1_INTERNAL_5 <= rfo2_data1(6);
RFO2_DATA1_INTERNAL_6 <= rfo2_data1(7);
RFO2_DATA1_INTERNAL_7 <= rfo2_data1(8);
RFO2_DATA1_INTERNAL_8 <= rfo2_data1(9);
RFO2_DATA1_INTERNAL_9 <= rfo2_data1(10);
RFO2_DATA1_INTERNAL_10 <= rfo2_data1(11);
RFO2_DATA1_INTERNAL_11 <= rfo2_data1(12);
RFO2_DATA1_INTERNAL_12 <= rfo2_data1(13);
RFO2_DATA1_INTERNAL_13 <= rfo2_data1(14);
RFO2_DATA1_INTERNAL_14 <= rfo2_data1(15);
RFO2_DATA1_INTERNAL_15 <= rfo2_data1(16);
RFO2_DATA1_INTERNAL_16 <= rfo2_data1(17);
RFO2_DATA1_INTERNAL_17 <= rfo2_data1(18);
RFO2_DATA1_INTERNAL_18 <= rfo2_data1(19);
RFO2_DATA1_INTERNAL_19 <= rfo2_data1(20);
RFO2_DATA1_INTERNAL_20 <= rfo2_data1(21);
RFO2_DATA1_INTERNAL_21 <= rfo2_data1(22);
RFO2_DATA1_INTERNAL_22 <= rfo2_data1(23);
RFO2_DATA1_INTERNAL_23 <= rfo2_data1(24);
RFO2_DATA1_INTERNAL_24 <= rfo2_data1(25);
RFO2_DATA1_INTERNAL_25 <= rfo2_data1(26);
RFO2_DATA1_INTERNAL_26 <= rfo2_data1(27);
RFO2_DATA1_INTERNAL_27 <= rfo2_data1(28);
RFO2_DATA1_INTERNAL_28 <= rfo2_data1(29);
RFO2_DATA1_INTERNAL_29 <= rfo2_data1(30);
RFO2_DATA1_INTERNAL_30 <= rfo2_data1(31);
RFO2_DATA2_INTERNAL <= rfo2_data2(0);
RFO2_DATA2_INTERNAL_0 <= rfo2_data2(1);
RFO2_DATA2_INTERNAL_1 <= rfo2_data2(2);
RFO2_DATA2_INTERNAL_2 <= rfo2_data2(3);
RFO2_DATA2_INTERNAL_3 <= rfo2_data2(4);
RFO2_DATA2_INTERNAL_4 <= rfo2_data2(5);
RFO2_DATA2_INTERNAL_5 <= rfo2_data2(6);
RFO2_DATA2_INTERNAL_6 <= rfo2_data2(7);
RFO2_DATA2_INTERNAL_7 <= rfo2_data2(8);
RFO2_DATA2_INTERNAL_8 <= rfo2_data2(9);
RFO2_DATA2_INTERNAL_9 <= rfo2_data2(10);
RFO2_DATA2_INTERNAL_10 <= rfo2_data2(11);
RFO2_DATA2_INTERNAL_11 <= rfo2_data2(12);
RFO2_DATA2_INTERNAL_12 <= rfo2_data2(13);
RFO2_DATA2_INTERNAL_13 <= rfo2_data2(14);
RFO2_DATA2_INTERNAL_14 <= rfo2_data2(15);
RFO2_DATA2_INTERNAL_15 <= rfo2_data2(16);
RFO2_DATA2_INTERNAL_16 <= rfo2_data2(17);
RFO2_DATA2_INTERNAL_17 <= rfo2_data2(18);
RFO2_DATA2_INTERNAL_18 <= rfo2_data2(19);
RFO2_DATA2_INTERNAL_19 <= rfo2_data2(20);
RFO2_DATA2_INTERNAL_20 <= rfo2_data2(21);
RFO2_DATA2_INTERNAL_21 <= rfo2_data2(22);
RFO2_DATA2_INTERNAL_22 <= rfo2_data2(23);
RFO2_DATA2_INTERNAL_23 <= rfo2_data2(24);
RFO2_DATA2_INTERNAL_24 <= rfo2_data2(25);
RFO2_DATA2_INTERNAL_25 <= rfo2_data2(26);
RFO2_DATA2_INTERNAL_26 <= rfo2_data2(27);
RFO2_DATA2_INTERNAL_27 <= rfo2_data2(28);
RFO2_DATA2_INTERNAL_28 <= rfo2_data2(29);
RFO2_DATA2_INTERNAL_29 <= rfo2_data2(30);
RFO2_DATA2_INTERNAL_30 <= rfo2_data2(31);
end beh;

